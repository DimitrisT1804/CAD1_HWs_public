// Generated netlist by CADI API on Date: 2025-10-09 17:35:40 //

module c1908 (N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88, N91, N94, N99, N104, N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899);
input N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88, N91, N94, N99, N104;
output N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899;

sg13g2_nor2_1 U210 (.A(n203), .B(n204), .Y(N2899));
sg13g2_xnor2_1 U211 (.A(n205), .B(n206), .Y(n204));
sg13g2_xor2_1 U212 (.A(n207), .B(n208), .X(n206));
sg13g2_nor2b_1 U213 (.A(n209), .B_N(N79), .Y(n207));
sg13g2_xor2_1 U214 (.A(n210), .B(n211), .X(N2892));
sg13g2_mux2_1 U215 (.A0(n212), .A1(n213), .S(n214), .X(n211));
sg13g2_nor2_1 U216 (.A(n215), .B(n216), .Y(n214));
sg13g2_xnor2_1 U217 (.A(n217), .B(n218), .Y(n216));
sg13g2_nor2_1 U218 (.A(N66), .B(n219), .Y(n213));
sg13g2_a21oi_1 U219 (.A1(N104), .A2(n220), .B1(n215), .Y(n212));
sg13g2_nor2_1 U220 (.A(n219), .B(N91), .Y(n215));
sg13g2_nand2_1 U221 (.A(n219), .B(n221), .Y(n210));
sg13g2_xor2_1 U222 (.A(n222), .B(n223), .X(N2891));
sg13g2_nor2_1 U223 (.A(n224), .B(N104), .Y(n223));
sg13g2_xor2_1 U224 (.A(n225), .B(n226), .X(n222));
sg13g2_nor2_1 U225 (.A(n227), .B(n228), .Y(n226));
sg13g2_o21ai_1 U226 (.A1(N63), .A2(n219), .B1(n229), .Y(n225));
sg13g2_inv_1 U227 (.A(n227), .Y(n229));
sg13g2_nor2_1 U228 (.A(n219), .B(N88), .Y(n227));
sg13g2_nor2_1 U229 (.A(n203), .B(n230), .Y(N2890));
sg13g2_xnor2_1 U230 (.A(n231), .B(n232), .Y(n230));
sg13g2_nor2_1 U231 (.A(n233), .B(n209), .Y(n232));
sg13g2_nor2_1 U232 (.A(n203), .B(n234), .Y(N2889));
sg13g2_xnor2_1 U233 (.A(n235), .B(n236), .Y(n234));
sg13g2_nor2b_1 U234 (.A(n209), .B_N(N85), .Y(n236));
sg13g2_nor2_1 U235 (.A(n203), .B(n237), .Y(N2888));
sg13g2_xnor2_1 U236 (.A(n238), .B(n239), .Y(n237));
sg13g2_nor2b_1 U237 (.A(n209), .B_N(N82), .Y(n239));
sg13g2_nor2_1 U238 (.A(n203), .B(n240), .Y(N2887));
sg13g2_xor2_1 U239 (.A(n241), .B(n242), .X(n240));
sg13g2_nor2b_1 U240 (.A(n209), .B_N(N76), .Y(n242));
sg13g2_nor2_1 U241 (.A(n203), .B(n243), .Y(N2886));
sg13g2_xor2_1 U242 (.A(n244), .B(n245), .X(n243));
sg13g2_nor2_1 U243 (.A(n246), .B(n209), .Y(n245));
sg13g2_or2_1 U244 (.A(n247), .B(n248), .X(n209));
sg13g2_nor2_1 U245 (.A(n219), .B(N99), .Y(n203));
sg13g2_nand4_1 U246 (.A(n247), .B(n249), .C(n250), .D(n219), .Y(N2811));
sg13g2_inv_1 U247 (.A(N104), .Y(n219));
sg13g2_nand3_1 U248 (.A(n251), .B(n252), .C(n253), .Y(n250));
sg13g2_a21oi_1 U249 (.A1(n254), .A2(n255), .B1(n256), .Y(n253));
sg13g2_o21ai_1 U250 (.A1(n257), .A2(n258), .B1(n259), .Y(n255));
sg13g2_o21ai_1 U251 (.A1(n260), .A2(n261), .B1(n262), .Y(n254));
sg13g2_nand3_1 U252 (.A(n262), .B(n263), .C(n259), .Y(n249));
sg13g2_o21ai_1 U253 (.A1(n256), .A2(n264), .B1(n265), .Y(n263));
sg13g2_o21ai_1 U254 (.A1(n266), .A2(n267), .B1(n251), .Y(n265));
sg13g2_inv_1 U255 (.A(n268), .Y(n251));
sg13g2_inv_1 U256 (.A(n269), .Y(n267));
sg13g2_o21ai_1 U257 (.A1(n270), .A2(n271), .B1(n272), .Y(n269));
sg13g2_a21oi_1 U258 (.A1(n273), .A2(n274), .B1(n264), .Y(n266));
sg13g2_inv_1 U259 (.A(n252), .Y(n264));
sg13g2_nor2b_1 U260 (.A(n221), .B_N(n224), .Y(n247));
sg13g2_nand2_1 U261 (.A(n275), .B(n276), .Y(n221));
sg13g2_and4_1 U262 (.A(n277), .B(n278), .C(n279), .D(n280), .X(n276));
sg13g2_and4_1 U263 (.A(n281), .B(n282), .C(n283), .D(n284), .X(n275));
sg13g2_and4_1 U264 (.A(n285), .B(n286), .C(n287), .D(n288), .X(n224));
sg13g2_and4_1 U265 (.A(n289), .B(n290), .C(n291), .D(n292), .X(n288));
sg13g2_and2_1 U266 (.A(n293), .B(n294), .X(n287));
sg13g2_xor2_1 U267 (.A(n295), .B(n284), .X(N2787));
sg13g2_nand3_1 U268 (.A(n296), .B(n297), .C(n252), .Y(n284));
sg13g2_xnor2_1 U269 (.A(N37), .B(n283), .Y(N2786));
sg13g2_nand3_1 U270 (.A(n298), .B(n262), .C(n252), .Y(n283));
sg13g2_xnor2_1 U271 (.A(N34), .B(n282), .Y(N2785));
sg13g2_nand3_1 U272 (.A(n299), .B(n257), .C(n252), .Y(n282));
sg13g2_xor2_1 U273 (.A(n300), .B(n281), .X(N2784));
sg13g2_nand3_1 U274 (.A(n299), .B(n258), .C(n252), .Y(n281));
sg13g2_a21oi_1 U275 (.A1(n301), .A2(N53), .B1(n302), .Y(n252));
sg13g2_xor2_1 U276 (.A(n303), .B(n280), .X(N2783));
sg13g2_nand4_1 U277 (.A(n296), .B(n272), .C(n271), .D(n304), .Y(n280));
sg13g2_inv_1 U278 (.A(n256), .Y(n272));
sg13g2_and3_1 U279 (.A(n261), .B(n305), .C(n258), .X(n296));
sg13g2_xnor2_1 U280 (.A(N22), .B(n292), .Y(N2782));
sg13g2_nand4_1 U281 (.A(n306), .B(n259), .C(n307), .D(n308), .Y(n292));
sg13g2_xnor2_1 U282 (.A(N19), .B(n291), .Y(N2781));
sg13g2_nand4_1 U283 (.A(n306), .B(n262), .C(n309), .D(n305), .Y(n291));
sg13g2_xnor2_1 U284 (.A(N16), .B(n290), .Y(N2780));
sg13g2_nand3_1 U285 (.A(n257), .B(n260), .C(n306), .Y(n290));
sg13g2_xnor2_1 U286 (.A(N13), .B(n289), .Y(N2779));
sg13g2_nand3_1 U287 (.A(n258), .B(n260), .C(n306), .Y(n289));
sg13g2_nor2b_1 U288 (.A(n256), .B_N(n310), .Y(n306));
sg13g2_nand2b_1 U289 (.A_N(n273), .B(n311), .Y(n256));
sg13g2_xnor2_1 U290 (.A(N46), .B(n279), .Y(N2768));
sg13g2_nand3_1 U291 (.A(n258), .B(n271), .C(n298), .Y(n279));
sg13g2_xnor2_1 U292 (.A(N43), .B(n278), .Y(N2767));
sg13g2_nand4_1 U293 (.A(n299), .B(n271), .C(n307), .D(n308), .Y(n278));
sg13g2_and2_1 U294 (.A(n297), .B(n260), .X(n299));
sg13g2_xnor2_1 U295 (.A(N28), .B(n277), .Y(N2762));
sg13g2_nand3_1 U296 (.A(n257), .B(n271), .C(n298), .Y(n277));
sg13g2_and3_1 U297 (.A(n309), .B(n305), .C(n297), .X(n298));
sg13g2_nor2b_1 U298 (.A(n274), .B_N(n304), .Y(n297));
sg13g2_o21ai_1 U299 (.A1(N91), .A2(n312), .B1(n268), .Y(n304));
sg13g2_xnor2_1 U300 (.A(N10), .B(n285), .Y(N2756));
sg13g2_nand4_1 U301 (.A(n261), .B(n262), .C(n313), .D(n305), .Y(n285));
sg13g2_xnor2_1 U302 (.A(N7), .B(n286), .Y(N2755));
sg13g2_nand3_1 U303 (.A(n259), .B(n313), .C(n257), .Y(n286));
sg13g2_nor2b_1 U304 (.A(n308), .B_N(n307), .Y(n257));
sg13g2_xnor2_1 U305 (.A(N4), .B(n294), .Y(N2754));
sg13g2_nand3_1 U306 (.A(n258), .B(n313), .C(n259), .Y(n294));
sg13g2_nor2_1 U307 (.A(n309), .B(n305), .Y(n259));
sg13g2_inv_1 U308 (.A(n261), .Y(n309));
sg13g2_nor2b_1 U309 (.A(n307), .B_N(n308), .Y(n258));
sg13g2_xnor2_1 U310 (.A(N1), .B(n293), .Y(N2753));
sg13g2_nand3_1 U311 (.A(n262), .B(n313), .C(n260), .Y(n293));
sg13g2_nor2_1 U312 (.A(n305), .B(n261), .Y(n260));
sg13g2_xnor2_1 U313 (.A(N79), .B(n314), .Y(n261));
sg13g2_nor2_1 U314 (.A(N94), .B(n315), .Y(n314));
sg13g2_xnor2_1 U315 (.A(n208), .B(n205), .Y(n315));
sg13g2_xnor2_1 U316 (.A(n316), .B(N1), .Y(n205));
sg13g2_nand2_1 U317 (.A(N49), .B(n317), .Y(n316));
sg13g2_xnor2_1 U318 (.A(n217), .B(n318), .Y(n208));
sg13g2_xor2_1 U319 (.A(n319), .B(n233), .X(n305));
sg13g2_o21ai_1 U320 (.A1(N94), .A2(n320), .B1(N56), .Y(n233));
sg13g2_nand2_1 U321 (.A(n231), .B(n248), .Y(n319));
sg13g2_xnor2_1 U322 (.A(n321), .B(n322), .Y(n231));
sg13g2_xor2_1 U323 (.A(N19), .B(n323), .X(n322));
sg13g2_xor2_1 U324 (.A(N37), .B(N28), .X(n323));
sg13g2_xor2_1 U325 (.A(n324), .B(n325), .X(n321));
sg13g2_xnor2_1 U326 (.A(N10), .B(n326), .Y(n325));
sg13g2_nand2_1 U327 (.A(N60), .B(n327), .Y(n326));
sg13g2_nor2b_1 U328 (.A(n274), .B_N(n310), .Y(n313));
sg13g2_nand2_1 U329 (.A(n273), .B(n311), .Y(n274));
sg13g2_o21ai_1 U330 (.A1(N94), .A2(n320), .B1(N60), .Y(n311));
sg13g2_xor2_1 U331 (.A(N76), .B(n328), .X(n273));
sg13g2_nor2_1 U332 (.A(N94), .B(n241), .Y(n328));
sg13g2_xor2_1 U333 (.A(n329), .B(n330), .X(n241));
sg13g2_xor2_1 U334 (.A(n331), .B(n332), .X(n330));
sg13g2_xor2_1 U335 (.A(N40), .B(N10), .X(n332));
sg13g2_nor2_1 U336 (.A(N104), .B(n220), .Y(n331));
sg13g2_inv_1 U337 (.A(N66), .Y(n220));
sg13g2_xor2_1 U338 (.A(n217), .B(n333), .X(n329));
sg13g2_xor2_1 U339 (.A(n334), .B(n335), .X(n217));
sg13g2_xor2_1 U340 (.A(N37), .B(N34), .X(n335));
sg13g2_xor2_1 U341 (.A(n336), .B(n300), .X(n334));
sg13g2_inv_1 U342 (.A(N31), .Y(n300));
sg13g2_and2_1 U343 (.A(n337), .B(n271), .X(n310));
sg13g2_a21oi_1 U344 (.A1(n301), .A2(N53), .B1(n270), .Y(n271));
sg13g2_inv_1 U345 (.A(n302), .Y(n270));
sg13g2_xnor2_1 U346 (.A(n246), .B(n338), .Y(n302));
sg13g2_nor2_1 U347 (.A(N94), .B(n244), .Y(n338));
sg13g2_xor2_1 U348 (.A(n339), .B(n340), .X(n244));
sg13g2_xor2_1 U349 (.A(N25), .B(n341), .X(n340));
sg13g2_nor2b_1 U350 (.A(N104), .B_N(N63), .Y(n341));
sg13g2_xnor2_1 U351 (.A(n228), .B(n336), .Y(n339));
sg13g2_xor2_1 U352 (.A(N28), .B(n342), .X(n336));
sg13g2_xor2_1 U353 (.A(N46), .B(N43), .X(n342));
sg13g2_xnor2_1 U354 (.A(n343), .B(n344), .Y(n228));
sg13g2_xor2_1 U355 (.A(N22), .B(N10), .X(n344));
sg13g2_xnor2_1 U356 (.A(n333), .B(n318), .Y(n343));
sg13g2_xor2_1 U357 (.A(N13), .B(n345), .X(n318));
sg13g2_xor2_1 U358 (.A(N19), .B(N16), .X(n345));
sg13g2_xor2_1 U359 (.A(N1), .B(n346), .X(n333));
sg13g2_xor2_1 U360 (.A(N7), .B(N4), .X(n346));
sg13g2_nand2_1 U361 (.A(n301), .B(N49), .Y(n246));
sg13g2_or2_1 U362 (.A(N72), .B(N94), .X(n301));
sg13g2_o21ai_1 U363 (.A1(N88), .A2(n312), .B1(n268), .Y(n337));
sg13g2_nand2_1 U364 (.A(n347), .B(N99), .Y(n268));
sg13g2_a21oi_1 U365 (.A1(N72), .A2(N69), .B1(N104), .Y(n347));
sg13g2_nand3_1 U366 (.A(N104), .B(n348), .C(N94), .Y(n312));
sg13g2_nand2_1 U367 (.A(N72), .B(N69), .Y(n348));
sg13g2_nor2_1 U368 (.A(n308), .B(n307), .Y(n262));
sg13g2_xnor2_1 U369 (.A(n349), .B(N85), .Y(n307));
sg13g2_nand2_1 U370 (.A(n235), .B(n248), .Y(n349));
sg13g2_xnor2_1 U371 (.A(n350), .B(n351), .Y(n235));
sg13g2_xor2_1 U372 (.A(n352), .B(n353), .X(n351));
sg13g2_xor2_1 U373 (.A(N34), .B(N28), .X(n353));
sg13g2_xor2_1 U374 (.A(N7), .B(N43), .X(n352));
sg13g2_xor2_1 U375 (.A(n354), .B(n355), .X(n350));
sg13g2_xor2_1 U376 (.A(N22), .B(N16), .X(n355));
sg13g2_nand2_1 U377 (.A(n327), .B(N56), .Y(n354));
sg13g2_nor2_1 U378 (.A(n320), .B(N104), .Y(n327));
sg13g2_inv_1 U379 (.A(N69), .Y(n320));
sg13g2_xnor2_1 U380 (.A(n356), .B(N82), .Y(n308));
sg13g2_nand2_1 U381 (.A(n238), .B(n248), .Y(n356));
sg13g2_inv_1 U382 (.A(N94), .Y(n248));
sg13g2_xnor2_1 U383 (.A(n357), .B(n358), .Y(n238));
sg13g2_xor2_1 U384 (.A(n359), .B(n360), .X(n358));
sg13g2_xor2_1 U385 (.A(N31), .B(N22), .X(n360));
sg13g2_xor2_1 U386 (.A(N43), .B(N4), .X(n359));
sg13g2_xor2_1 U387 (.A(n324), .B(n361), .X(n357));
sg13g2_xnor2_1 U388 (.A(N13), .B(n362), .Y(n361));
sg13g2_nand2_1 U389 (.A(N53), .B(n317), .Y(n362));
sg13g2_nor2_1 U390 (.A(N104), .B(N72), .Y(n317));
sg13g2_xnor2_1 U391 (.A(N46), .B(n218), .Y(n324));
sg13g2_xor2_1 U392 (.A(n303), .B(n295), .X(n218));
sg13g2_inv_1 U393 (.A(N40), .Y(n295));
sg13g2_inv_1 U394 (.A(N25), .Y(n303));
endmodule

