// Generated netlist by CADI API on Date: 2025-10-16 19:07:31 //

module aes192 (clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_i_8_, data_i_9_, data_i_10_, data_i_11_, data_i_12_, data_i_13_, data_i_14_, data_i_15_, data_i_16_, data_i_17_, data_i_18_, data_i_19_, data_i_20_, data_i_21_, data_i_22_, data_i_23_, data_i_24_, data_i_25_, data_i_26_, data_i_27_, data_i_28_, data_i_29_, data_i_30_, data_i_31_, data_i_32_, data_i_33_, data_i_34_, data_i_35_, data_i_36_, data_i_37_, data_i_38_, data_i_39_, data_i_40_, data_i_41_, data_i_42_, data_i_43_, data_i_44_, data_i_45_, data_i_46_, data_i_47_, data_i_48_, data_i_49_, data_i_50_, data_i_51_, data_i_52_, data_i_53_, data_i_54_, data_i_55_, data_i_56_, data_i_57_, data_i_58_, data_i_59_, data_i_60_, data_i_61_, data_i_62_, data_i_63_, data_i_64_, data_i_65_, data_i_66_, data_i_67_, data_i_68_, data_i_69_, data_i_70_, data_i_71_, data_i_72_, data_i_73_, data_i_74_, data_i_75_, data_i_76_, data_i_77_, data_i_78_, data_i_79_, data_i_80_, data_i_81_, data_i_82_, data_i_83_, data_i_84_, data_i_85_, data_i_86_, data_i_87_, data_i_88_, data_i_89_, data_i_90_, data_i_91_, data_i_92_, data_i_93_, data_i_94_, data_i_95_, data_i_96_, data_i_97_, data_i_98_, data_i_99_, data_i_100_, data_i_101_, data_i_102_, data_i_103_, data_i_104_, data_i_105_, data_i_106_, data_i_107_, data_i_108_, data_i_109_, data_i_110_, data_i_111_, data_i_112_, data_i_113_, data_i_114_, data_i_115_, data_i_116_, data_i_117_, data_i_118_, data_i_119_, data_i_120_, data_i_121_, data_i_122_, data_i_123_, data_i_124_, data_i_125_, data_i_126_, data_i_127_, data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_, data_o_32_, data_o_33_, data_o_34_, data_o_35_, data_o_36_, data_o_37_, data_o_38_, data_o_39_, data_o_40_, data_o_41_, data_o_42_, data_o_43_, data_o_44_, data_o_45_, data_o_46_, data_o_47_, data_o_48_, data_o_49_, data_o_50_, data_o_51_, data_o_52_, data_o_53_, data_o_54_, data_o_55_, data_o_56_, data_o_57_, data_o_58_, data_o_59_, data_o_60_, data_o_61_, data_o_62_, data_o_63_, data_o_64_, data_o_65_, data_o_66_, data_o_67_, data_o_68_, data_o_69_, data_o_70_, data_o_71_, data_o_72_, data_o_73_, data_o_74_, data_o_75_, data_o_76_, data_o_77_, data_o_78_, data_o_79_, data_o_80_, data_o_81_, data_o_82_, data_o_83_, data_o_84_, data_o_85_, data_o_86_, data_o_87_, data_o_88_, data_o_89_, data_o_90_, data_o_91_, data_o_92_, data_o_93_, data_o_94_, data_o_95_, data_o_96_, data_o_97_, data_o_98_, data_o_99_, data_o_100_, data_o_101_, data_o_102_, data_o_103_, data_o_104_, data_o_105_, data_o_106_, data_o_107_, data_o_108_, data_o_109_, data_o_110_, data_o_111_, data_o_112_, data_o_113_, data_o_114_, data_o_115_, data_o_116_, data_o_117_, data_o_118_, data_o_119_, data_o_120_, data_o_121_, data_o_122_, data_o_123_, data_o_124_, data_o_125_, data_o_126_, data_o_127_, decrypt_i, key_i_0_, key_i_1_, key_i_2_, key_i_3_, key_i_4_, key_i_5_, key_i_6_, key_i_7_, key_i_8_, key_i_9_, key_i_10_, key_i_11_, key_i_12_, key_i_13_, key_i_14_, key_i_15_, key_i_16_, key_i_17_, key_i_18_, key_i_19_, key_i_20_, key_i_21_, key_i_22_, key_i_23_, key_i_24_, key_i_25_, key_i_26_, key_i_27_, key_i_28_, key_i_29_, key_i_30_, key_i_31_, key_i_32_, key_i_33_, key_i_34_, key_i_35_, key_i_36_, key_i_37_, key_i_38_, key_i_39_, key_i_40_, key_i_41_, key_i_42_, key_i_43_, key_i_44_, key_i_45_, key_i_46_, key_i_47_, key_i_48_, key_i_49_, key_i_50_, key_i_51_, key_i_52_, key_i_53_, key_i_54_, key_i_55_, key_i_56_, key_i_57_, key_i_58_, key_i_59_, key_i_60_, key_i_61_, key_i_62_, key_i_63_, key_i_64_, key_i_65_, key_i_66_, key_i_67_, key_i_68_, key_i_69_, key_i_70_, key_i_71_, key_i_72_, key_i_73_, key_i_74_, key_i_75_, key_i_76_, key_i_77_, key_i_78_, key_i_79_, key_i_80_, key_i_81_, key_i_82_, key_i_83_, key_i_84_, key_i_85_, key_i_86_, key_i_87_, key_i_88_, key_i_89_, key_i_90_, key_i_91_, key_i_92_, key_i_93_, key_i_94_, key_i_95_, key_i_96_, key_i_97_, key_i_98_, key_i_99_, key_i_100_, key_i_101_, key_i_102_, key_i_103_, key_i_104_, key_i_105_, key_i_106_, key_i_107_, key_i_108_, key_i_109_, key_i_110_, key_i_111_, key_i_112_, key_i_113_, key_i_114_, key_i_115_, key_i_116_, key_i_117_, key_i_118_, key_i_119_, key_i_120_, key_i_121_, key_i_122_, key_i_123_, key_i_124_, key_i_125_, key_i_126_, key_i_127_, key_i_128_, key_i_129_, key_i_130_, key_i_131_, key_i_132_, key_i_133_, key_i_134_, key_i_135_, key_i_136_, key_i_137_, key_i_138_, key_i_139_, key_i_140_, key_i_141_, key_i_142_, key_i_143_, key_i_144_, key_i_145_, key_i_146_, key_i_147_, key_i_148_, key_i_149_, key_i_150_, key_i_151_, key_i_152_, key_i_153_, key_i_154_, key_i_155_, key_i_156_, key_i_157_, key_i_158_, key_i_159_, key_i_160_, key_i_161_, key_i_162_, key_i_163_, key_i_164_, key_i_165_, key_i_166_, key_i_167_, key_i_168_, key_i_169_, key_i_170_, key_i_171_, key_i_172_, key_i_173_, key_i_174_, key_i_175_, key_i_176_, key_i_177_, key_i_178_, key_i_179_, key_i_180_, key_i_181_, key_i_182_, key_i_183_, key_i_184_, key_i_185_, key_i_186_, key_i_187_, key_i_188_, key_i_189_, key_i_190_, key_i_191_, load_i, ready_o, reset);
input clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_i_8_, data_i_9_, data_i_10_, data_i_11_, data_i_12_, data_i_13_, data_i_14_, data_i_15_, data_i_16_, data_i_17_, data_i_18_, data_i_19_, data_i_20_, data_i_21_, data_i_22_, data_i_23_, data_i_24_, data_i_25_, data_i_26_, data_i_27_, data_i_28_, data_i_29_, data_i_30_, data_i_31_, data_i_32_, data_i_33_, data_i_34_, data_i_35_, data_i_36_, data_i_37_, data_i_38_, data_i_39_, data_i_40_, data_i_41_, data_i_42_, data_i_43_, data_i_44_, data_i_45_, data_i_46_, data_i_47_, data_i_48_, data_i_49_, data_i_50_, data_i_51_, data_i_52_, data_i_53_, data_i_54_, data_i_55_, data_i_56_, data_i_57_, data_i_58_, data_i_59_, data_i_60_, data_i_61_, data_i_62_, data_i_63_, data_i_64_, data_i_65_, data_i_66_, data_i_67_, data_i_68_, data_i_69_, data_i_70_, data_i_71_, data_i_72_, data_i_73_, data_i_74_, data_i_75_, data_i_76_, data_i_77_, data_i_78_, data_i_79_, data_i_80_, data_i_81_, data_i_82_, data_i_83_, data_i_84_, data_i_85_, data_i_86_, data_i_87_, data_i_88_, data_i_89_, data_i_90_, data_i_91_, data_i_92_, data_i_93_, data_i_94_, data_i_95_, data_i_96_, data_i_97_, data_i_98_, data_i_99_, data_i_100_, data_i_101_, data_i_102_, data_i_103_, data_i_104_, data_i_105_, data_i_106_, data_i_107_, data_i_108_, data_i_109_, data_i_110_, data_i_111_, data_i_112_, data_i_113_, data_i_114_, data_i_115_, data_i_116_, data_i_117_, data_i_118_, data_i_119_, data_i_120_, data_i_121_, data_i_122_, data_i_123_, data_i_124_, data_i_125_, data_i_126_, data_i_127_, decrypt_i, key_i_0_, key_i_1_, key_i_2_, key_i_3_, key_i_4_, key_i_5_, key_i_6_, key_i_7_, key_i_8_, key_i_9_, key_i_10_, key_i_11_, key_i_12_, key_i_13_, key_i_14_, key_i_15_, key_i_16_, key_i_17_, key_i_18_, key_i_19_, key_i_20_, key_i_21_, key_i_22_, key_i_23_, key_i_24_, key_i_25_, key_i_26_, key_i_27_, key_i_28_, key_i_29_, key_i_30_, key_i_31_, key_i_32_, key_i_33_, key_i_34_, key_i_35_, key_i_36_, key_i_37_, key_i_38_, key_i_39_, key_i_40_, key_i_41_, key_i_42_, key_i_43_, key_i_44_, key_i_45_, key_i_46_, key_i_47_, key_i_48_, key_i_49_, key_i_50_, key_i_51_, key_i_52_, key_i_53_, key_i_54_, key_i_55_, key_i_56_, key_i_57_, key_i_58_, key_i_59_, key_i_60_, key_i_61_, key_i_62_, key_i_63_, key_i_64_, key_i_65_, key_i_66_, key_i_67_, key_i_68_, key_i_69_, key_i_70_, key_i_71_, key_i_72_, key_i_73_, key_i_74_, key_i_75_, key_i_76_, key_i_77_, key_i_78_, key_i_79_, key_i_80_, key_i_81_, key_i_82_, key_i_83_, key_i_84_, key_i_85_, key_i_86_, key_i_87_, key_i_88_, key_i_89_, key_i_90_, key_i_91_, key_i_92_, key_i_93_, key_i_94_, key_i_95_, key_i_96_, key_i_97_, key_i_98_, key_i_99_, key_i_100_, key_i_101_, key_i_102_, key_i_103_, key_i_104_, key_i_105_, key_i_106_, key_i_107_, key_i_108_, key_i_109_, key_i_110_, key_i_111_, key_i_112_, key_i_113_, key_i_114_, key_i_115_, key_i_116_, key_i_117_, key_i_118_, key_i_119_, key_i_120_, key_i_121_, key_i_122_, key_i_123_, key_i_124_, key_i_125_, key_i_126_, key_i_127_, key_i_128_, key_i_129_, key_i_130_, key_i_131_, key_i_132_, key_i_133_, key_i_134_, key_i_135_, key_i_136_, key_i_137_, key_i_138_, key_i_139_, key_i_140_, key_i_141_, key_i_142_, key_i_143_, key_i_144_, key_i_145_, key_i_146_, key_i_147_, key_i_148_, key_i_149_, key_i_150_, key_i_151_, key_i_152_, key_i_153_, key_i_154_, key_i_155_, key_i_156_, key_i_157_, key_i_158_, key_i_159_, key_i_160_, key_i_161_, key_i_162_, key_i_163_, key_i_164_, key_i_165_, key_i_166_, key_i_167_, key_i_168_, key_i_169_, key_i_170_, key_i_171_, key_i_172_, key_i_173_, key_i_174_, key_i_175_, key_i_176_, key_i_177_, key_i_178_, key_i_179_, key_i_180_, key_i_181_, key_i_182_, key_i_183_, key_i_184_, key_i_185_, key_i_186_, key_i_187_, key_i_188_, key_i_189_, key_i_190_, key_i_191_, load_i, reset;
output data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_, data_o_32_, data_o_33_, data_o_34_, data_o_35_, data_o_36_, data_o_37_, data_o_38_, data_o_39_, data_o_40_, data_o_41_, data_o_42_, data_o_43_, data_o_44_, data_o_45_, data_o_46_, data_o_47_, data_o_48_, data_o_49_, data_o_50_, data_o_51_, data_o_52_, data_o_53_, data_o_54_, data_o_55_, data_o_56_, data_o_57_, data_o_58_, data_o_59_, data_o_60_, data_o_61_, data_o_62_, data_o_63_, data_o_64_, data_o_65_, data_o_66_, data_o_67_, data_o_68_, data_o_69_, data_o_70_, data_o_71_, data_o_72_, data_o_73_, data_o_74_, data_o_75_, data_o_76_, data_o_77_, data_o_78_, data_o_79_, data_o_80_, data_o_81_, data_o_82_, data_o_83_, data_o_84_, data_o_85_, data_o_86_, data_o_87_, data_o_88_, data_o_89_, data_o_90_, data_o_91_, data_o_92_, data_o_93_, data_o_94_, data_o_95_, data_o_96_, data_o_97_, data_o_98_, data_o_99_, data_o_100_, data_o_101_, data_o_102_, data_o_103_, data_o_104_, data_o_105_, data_o_106_, data_o_107_, data_o_108_, data_o_109_, data_o_110_, data_o_111_, data_o_112_, data_o_113_, data_o_114_, data_o_115_, data_o_116_, data_o_117_, data_o_118_, data_o_119_, data_o_120_, data_o_121_, data_o_122_, data_o_123_, data_o_124_, data_o_125_, data_o_126_, data_o_127_, ready_o;

sg13g2_nand2_2 C3810 (.A(n3681), .B(N1628), .Y(n3695));
sg13g2_nand2_2 C3811 (.A(N1622), .B(N1625), .Y(n3696));
sg13g2_nand2_2 C3814 (.A(N1622), .B(N1628), .Y(n3699));
sg13g2_nand2_2 C3815 (.A(N1623), .B(N1625), .Y(n3700));
sg13g2_nand2_2 C3818 (.A(N1623), .B(N1628), .Y(n3732));
sg13g2_nand2_2 C3819 (.A(n3683), .B(N1625), .Y(n3703));
sg13g2_nand2_2 C3821 (.A(n3683), .B(N1627), .Y(n3731));
sg13g2_nand2_2 C3867 (.A(subbytes_ready_o), .B(N29), .Y(n3707));
sg13g2_nand2_2 C3871 (.A(mixcol_ready_o), .B(decrypt_i), .Y(n3710));
sg13g2_nand2_2 C3887 (.A(N29), .B(mixcol_ready_o), .Y(n554));
sg13g2_nand2_2 C3905 (.A(n3714), .B(n3715), .Y(N587));
sg13g2_nand2_2 C3906 (.A(N1594), .B(N29), .Y(n3714));
sg13g2_nand2_2 C3907 (.A(N1617), .B(decrypt_i), .Y(n3715));
sg13g2_nand2_2 C4300 (.A(N1617), .B(addroundkey_start_i), .Y(net24695));
sg13g2_nand2_2 C4301 (.A(addroundkey_start_i), .B(N1620), .Y(n168));
sg13g2_nand2_2 C4303 (.A(n3716), .B(n3721), .Y(N1645));
sg13g2_nand2_2 C4305 (.A(n3718), .B(n3719), .Y(N1641));
sg13g2_nand2_2 C4309 (.A(N1325), .B(N1125), .Y(n3721));
sg13g2_nand2_2 C4310 (.A(N1652), .B(keysched_ready_o), .Y(n166));
sg13g2_nand2_2 C4311 (.A(n3722), .B(n3727), .Y(N1652));
sg13g2_nand2_2 C4313 (.A(n4232), .B(n3725), .Y(N1648));
sg13g2_nand2_2 C4317 (.A(N1325), .B(N1124), .Y(n3727));
sg13g2_nand2_2 C4319 (.A(n3728), .B(n3734), .Y(N1659));
sg13g2_nand2_2 C4321 (.A(N1653), .B(N1654), .Y(n3729));
sg13g2_nand2_2 C4323 (.A(n3731), .B(n3732), .Y(N1654));
sg13g2_inv_4 I_7 (.A(N1589), .Y(N1590));
sg13g2_a21oi_1 U1 (.A1(n1), .A2(N1324), .B1(N1641), .Y(n3716));
sg13g2_nand3_1 U2 (.A(n1771), .B(n2), .C(n1770), .Y(next_addroundkey_data_reg_0));
sg13g2_nand3_1 U3 (.A(n1766), .B(n3), .C(n1765), .Y(next_addroundkey_data_reg_100));
sg13g2_nand3_1 U4 (.A(n1761), .B(n4), .C(n1760), .Y(next_addroundkey_data_reg_101));
sg13g2_nand3_1 U5 (.A(n1756), .B(n5), .C(n1755), .Y(next_addroundkey_data_reg_102));
sg13g2_nand3_1 U6 (.A(n1751), .B(n6), .C(n1750), .Y(next_addroundkey_data_reg_103));
sg13g2_nand3_1 U7 (.A(n1746), .B(n7), .C(n1745), .Y(next_addroundkey_data_reg_104));
sg13g2_nand3_1 U8 (.A(n1741), .B(n8), .C(n1740), .Y(next_addroundkey_data_reg_105));
sg13g2_o21ai_1 U9 (.A1(n4328), .A2(n558), .B1(n559), .Y(subbytes_data_i_9));
sg13g2_nand3_1 U10 (.A(n1736), .B(n9), .C(n1735), .Y(next_addroundkey_data_reg_106));
sg13g2_o21ai_1 U11 (.A1(n4327), .A2(n561), .B1(n562), .Y(subbytes_data_i_99));
sg13g2_nand2_2 U12 (.A(data_o_99_), .B(n4323), .Y(n562));
sg13g2_o21ai_1 U13 (.A1(n4325), .A2(n563), .B1(n564), .Y(subbytes_data_i_98));
sg13g2_nand2_2 U14 (.A(data_o_98_), .B(n4318), .Y(n564));
sg13g2_o21ai_1 U15 (.A1(n4326), .A2(n565), .B1(n566), .Y(subbytes_data_i_97));
sg13g2_nand2_2 U16 (.A(data_o_97_), .B(n4321), .Y(n566));
sg13g2_o21ai_1 U17 (.A1(n4325), .A2(n567), .B1(n568), .Y(subbytes_data_i_96));
sg13g2_nand2_2 U18 (.A(data_o_96_), .B(n4298), .Y(n568));
sg13g2_o21ai_1 U19 (.A1(n4328), .A2(n569), .B1(n570), .Y(subbytes_data_i_95));
sg13g2_nand2_2 U20 (.A(data_o_95_), .B(n4318), .Y(n570));
sg13g2_nand3_1 U21 (.A(n1731), .B(n10), .C(n1730), .Y(next_addroundkey_data_reg_107));
sg13g2_nand2_2 U22 (.A(data_o_94_), .B(n4323), .Y(n572));
sg13g2_nand3_1 U23 (.A(n1726), .B(n11), .C(n1725), .Y(next_addroundkey_data_reg_108));
sg13g2_nand2_2 U24 (.A(data_o_93_), .B(n4317), .Y(n574));
sg13g2_nand3_1 U25 (.A(n1721), .B(n12), .C(n1720), .Y(next_addroundkey_data_reg_109));
sg13g2_nand3_1 U26 (.A(n1716), .B(n13), .C(n1715), .Y(next_addroundkey_data_reg_10));
sg13g2_o21ai_1 U27 (.A1(n4329), .A2(n577), .B1(n578), .Y(subbytes_data_i_91));
sg13g2_nand3_1 U28 (.A(n1711), .B(n14), .C(n1710), .Y(next_addroundkey_data_reg_110));
sg13g2_o21ai_1 U29 (.A1(n4328), .A2(n579), .B1(n580), .Y(subbytes_data_i_90));
sg13g2_nand2_2 U30 (.A(data_o_90_), .B(n4319), .Y(n580));
sg13g2_o21ai_1 U31 (.A1(n4329), .A2(n581), .B1(n582), .Y(subbytes_data_i_8));
sg13g2_nand3_1 U32 (.A(n1706), .B(n15), .C(n1705), .Y(next_addroundkey_data_reg_111));
sg13g2_o21ai_1 U33 (.A1(n4329), .A2(n583), .B1(n584), .Y(subbytes_data_i_89));
sg13g2_nand2_2 U34 (.A(data_o_89_), .B(n4318), .Y(n584));
sg13g2_nand3_1 U35 (.A(n1701), .B(n16), .C(n1700), .Y(next_addroundkey_data_reg_112));
sg13g2_nand3_1 U36 (.A(n1696), .B(n17), .C(n1695), .Y(next_addroundkey_data_reg_113));
sg13g2_o21ai_1 U37 (.A1(n4327), .A2(n587), .B1(n588), .Y(subbytes_data_i_87));
sg13g2_nand2_2 U38 (.A(data_o_87_), .B(n4318), .Y(n588));
sg13g2_o21ai_1 U39 (.A1(n4327), .A2(n589), .B1(n590), .Y(subbytes_data_i_86));
sg13g2_nand3_1 U40 (.A(n1691), .B(n18), .C(n1690), .Y(next_addroundkey_data_reg_114));
sg13g2_nand3_1 U41 (.A(n1686), .B(n19), .C(n1685), .Y(next_addroundkey_data_reg_115));
sg13g2_nand3_1 U42 (.A(n1681), .B(n20), .C(n1680), .Y(next_addroundkey_data_reg_116));
sg13g2_o21ai_1 U43 (.A1(n4329), .A2(n593), .B1(n594), .Y(subbytes_data_i_84));
sg13g2_nand3_1 U44 (.A(n1676), .B(n21), .C(n1675), .Y(next_addroundkey_data_reg_117));
sg13g2_nand3_1 U45 (.A(n1671), .B(n22), .C(n1670), .Y(next_addroundkey_data_reg_118));
sg13g2_nand3_1 U46 (.A(n1666), .B(n23), .C(n1665), .Y(next_addroundkey_data_reg_119));
sg13g2_o21ai_1 U47 (.A1(n4328), .A2(n597), .B1(n598), .Y(subbytes_data_i_82));
sg13g2_nand3_1 U48 (.A(n1661), .B(n24), .C(n1660), .Y(next_addroundkey_data_reg_11));
sg13g2_o21ai_1 U49 (.A1(n4325), .A2(n599), .B1(n600), .Y(subbytes_data_i_81));
sg13g2_nand2_2 U50 (.A(data_o_81_), .B(n4318), .Y(n600));
sg13g2_o21ai_1 U51 (.A1(n4325), .A2(n601), .B1(n602), .Y(subbytes_data_i_80));
sg13g2_nand2_2 U52 (.A(data_o_80_), .B(n4320), .Y(n602));
sg13g2_o21ai_1 U53 (.A1(n4325), .A2(n603), .B1(n604), .Y(subbytes_data_i_7));
sg13g2_nand2_2 U54 (.A(data_o_7_), .B(n4323), .Y(n604));
sg13g2_nand3_1 U55 (.A(n1656), .B(n25), .C(n1655), .Y(next_addroundkey_data_reg_120));
sg13g2_nand2_2 U56 (.A(data_o_79_), .B(n4319), .Y(n606));
sg13g2_o21ai_1 U57 (.A1(n4325), .A2(n607), .B1(n608), .Y(subbytes_data_i_78));
sg13g2_nand3_1 U58 (.A(n1651), .B(n26), .C(n1650), .Y(next_addroundkey_data_reg_121));
sg13g2_nand3_1 U59 (.A(n1646), .B(n27), .C(n1645), .Y(next_addroundkey_data_reg_122));
sg13g2_nand3_1 U60 (.A(n1641), .B(n28), .C(n1640), .Y(next_addroundkey_data_reg_123));
sg13g2_nand3_1 U61 (.A(n1636), .B(n29), .C(n1635), .Y(next_addroundkey_data_reg_124));
sg13g2_nand3_1 U62 (.A(n1631), .B(n30), .C(n1630), .Y(next_addroundkey_data_reg_125));
sg13g2_nand3_1 U63 (.A(n1626), .B(n31), .C(n1625), .Y(next_addroundkey_data_reg_126));
sg13g2_nand2_2 U64 (.A(data_o_75_), .B(n4317), .Y(n614));
sg13g2_o21ai_1 U65 (.A1(n4325), .A2(n615), .B1(n616), .Y(subbytes_data_i_74));
sg13g2_nand2_2 U66 (.A(data_o_74_), .B(n4319), .Y(n616));
sg13g2_nand3_1 U67 (.A(n1621), .B(n32), .C(n1620), .Y(next_addroundkey_data_reg_127));
sg13g2_nand2_2 U68 (.A(data_o_73_), .B(n4318), .Y(n618));
sg13g2_nand3_1 U69 (.A(n1616), .B(n33), .C(n1615), .Y(next_addroundkey_data_reg_12));
sg13g2_nand3_1 U70 (.A(n1611), .B(n34), .C(n1610), .Y(next_addroundkey_data_reg_13));
sg13g2_o21ai_1 U71 (.A1(n4325), .A2(n621), .B1(n622), .Y(subbytes_data_i_71));
sg13g2_nand2_2 U72 (.A(data_o_71_), .B(n4317), .Y(n622));
sg13g2_o21ai_1 U73 (.A1(n4325), .A2(n623), .B1(n624), .Y(subbytes_data_i_70));
sg13g2_nand2_2 U74 (.A(data_o_70_), .B(n4298), .Y(n624));
sg13g2_o21ai_1 U75 (.A1(n4327), .A2(n625), .B1(n626), .Y(subbytes_data_i_6));
sg13g2_nand3_1 U76 (.A(n1606), .B(n35), .C(n1605), .Y(next_addroundkey_data_reg_14));
sg13g2_nand3_1 U77 (.A(n1601), .B(n36), .C(n1600), .Y(next_addroundkey_data_reg_15));
sg13g2_nand3_1 U78 (.A(n1596), .B(n165), .C(n1595), .Y(next_addroundkey_data_reg_16));
sg13g2_nand3_1 U79 (.A(n1591), .B(n167), .C(n1590), .Y(next_addroundkey_data_reg_17));
sg13g2_nand3_1 U80 (.A(n1586), .B(n435), .C(n1585), .Y(next_addroundkey_data_reg_18));
sg13g2_o21ai_1 U81 (.A1(n4326), .A2(n631), .B1(n632), .Y(subbytes_data_i_67));
sg13g2_nand2_2 U82 (.A(data_o_67_), .B(n4321), .Y(n632));
sg13g2_o21ai_1 U83 (.A1(n4325), .A2(n633), .B1(n634), .Y(subbytes_data_i_66));
sg13g2_nand2_2 U84 (.A(data_o_66_), .B(n4319), .Y(n634));
sg13g2_nand3_1 U85 (.A(n1581), .B(n436), .C(n1580), .Y(next_addroundkey_data_reg_19));
sg13g2_nand2_2 U86 (.A(data_o_65_), .B(n4323), .Y(n636));
sg13g2_nand3_1 U87 (.A(n1576), .B(n529), .C(n1575), .Y(next_addroundkey_data_reg_1));
sg13g2_nand3_1 U88 (.A(n1571), .B(n530), .C(n1570), .Y(next_addroundkey_data_reg_20));
sg13g2_nand3_1 U89 (.A(n1566), .B(n531), .C(n1565), .Y(next_addroundkey_data_reg_21));
sg13g2_nand3_1 U90 (.A(n1561), .B(n532), .C(n1560), .Y(next_addroundkey_data_reg_22));
sg13g2_o21ai_1 U91 (.A1(n4330), .A2(n641), .B1(n642), .Y(subbytes_data_i_62));
sg13g2_nand2_2 U92 (.A(data_o_62_), .B(n4323), .Y(n642));
sg13g2_o21ai_1 U93 (.A1(n4328), .A2(n643), .B1(n644), .Y(subbytes_data_i_61));
sg13g2_nand2_2 U94 (.A(data_o_61_), .B(n4323), .Y(n644));
sg13g2_nand3_1 U95 (.A(n1556), .B(n533), .C(n1555), .Y(next_addroundkey_data_reg_23));
sg13g2_nand2_2 U96 (.A(data_o_60_), .B(n4316), .Y(n646));
sg13g2_o21ai_1 U97 (.A1(n4326), .A2(n647), .B1(n648), .Y(subbytes_data_i_5));
sg13g2_nand2_2 U98 (.A(data_o_5_), .B(n4320), .Y(n648));
sg13g2_o21ai_1 U99 (.A1(n4326), .A2(n649), .B1(n650), .Y(subbytes_data_i_59));
sg13g2_nand3_1 U100 (.A(n1551), .B(n534), .C(n1550), .Y(next_addroundkey_data_reg_24));
sg13g2_o21ai_1 U101 (.A1(n4326), .A2(n651), .B1(n652), .Y(subbytes_data_i_58));
sg13g2_nand2_2 U102 (.A(data_o_58_), .B(n4318), .Y(n652));
sg13g2_o21ai_1 U103 (.A1(n4326), .A2(n653), .B1(n654), .Y(subbytes_data_i_57));
sg13g2_nand2_2 U104 (.A(data_o_57_), .B(n4319), .Y(n654));
sg13g2_o21ai_1 U105 (.A1(n4326), .A2(n655), .B1(n656), .Y(subbytes_data_i_56));
sg13g2_nand2_2 U106 (.A(data_o_56_), .B(n4321), .Y(n656));
sg13g2_nand3_1 U107 (.A(n1546), .B(n535), .C(n1545), .Y(next_addroundkey_data_reg_25));
sg13g2_nand2_2 U108 (.A(data_o_55_), .B(n4298), .Y(n658));
sg13g2_o21ai_1 U109 (.A1(n4326), .A2(n659), .B1(n660), .Y(subbytes_data_i_54));
sg13g2_nand2_2 U110 (.A(data_o_54_), .B(n4321), .Y(n660));
sg13g2_o21ai_1 U111 (.A1(n4326), .A2(n661), .B1(n662), .Y(subbytes_data_i_53));
sg13g2_nand2_2 U112 (.A(data_o_53_), .B(n4319), .Y(n662));
sg13g2_o21ai_1 U113 (.A1(n4326), .A2(n663), .B1(n664), .Y(subbytes_data_i_52));
sg13g2_nand2_2 U114 (.A(data_o_52_), .B(n4298), .Y(n664));
sg13g2_o21ai_1 U115 (.A1(n4326), .A2(n665), .B1(n666), .Y(subbytes_data_i_51));
sg13g2_nand2_2 U116 (.A(data_o_51_), .B(n4320), .Y(n666));
sg13g2_o21ai_1 U117 (.A1(n4326), .A2(n667), .B1(n668), .Y(subbytes_data_i_50));
sg13g2_nand2_2 U118 (.A(data_o_50_), .B(n4319), .Y(n668));
sg13g2_o21ai_1 U119 (.A1(n4327), .A2(n669), .B1(n670), .Y(subbytes_data_i_4));
sg13g2_nand2_2 U120 (.A(data_o_4_), .B(n4298), .Y(n670));
sg13g2_o21ai_1 U121 (.A1(n4329), .A2(n671), .B1(n672), .Y(subbytes_data_i_49));
sg13g2_nand2_2 U122 (.A(data_o_49_), .B(n4319), .Y(n672));
sg13g2_o21ai_1 U123 (.A1(n4328), .A2(n673), .B1(n674), .Y(subbytes_data_i_48));
sg13g2_nand3_1 U124 (.A(n1541), .B(n536), .C(n1540), .Y(next_addroundkey_data_reg_26));
sg13g2_nand3_1 U125 (.A(n1536), .B(n537), .C(n1535), .Y(next_addroundkey_data_reg_27));
sg13g2_nand3_1 U126 (.A(n1531), .B(n538), .C(n1530), .Y(next_addroundkey_data_reg_28));
sg13g2_o21ai_1 U127 (.A1(n4326), .A2(n677), .B1(n678), .Y(subbytes_data_i_46));
sg13g2_nand2_2 U128 (.A(data_o_46_), .B(n4298), .Y(n678));
sg13g2_o21ai_1 U129 (.A1(n4328), .A2(n679), .B1(n680), .Y(subbytes_data_i_45));
sg13g2_nand2_2 U130 (.A(data_o_45_), .B(n4298), .Y(n680));
sg13g2_o21ai_1 U131 (.A1(n4329), .A2(n681), .B1(n682), .Y(subbytes_data_i_44));
sg13g2_nand2_2 U132 (.A(data_o_44_), .B(n4321), .Y(n682));
sg13g2_o21ai_1 U133 (.A1(n4325), .A2(n683), .B1(n684), .Y(subbytes_data_i_43));
sg13g2_nand2_2 U134 (.A(data_o_43_), .B(n4298), .Y(n684));
sg13g2_o21ai_1 U135 (.A1(n4330), .A2(n685), .B1(n686), .Y(subbytes_data_i_42));
sg13g2_nand2_2 U136 (.A(data_o_42_), .B(n4321), .Y(n686));
sg13g2_o21ai_1 U137 (.A1(n4326), .A2(n687), .B1(n688), .Y(subbytes_data_i_41));
sg13g2_nand2_2 U138 (.A(data_o_41_), .B(n4321), .Y(n688));
sg13g2_o21ai_1 U139 (.A1(n4326), .A2(n689), .B1(n690), .Y(subbytes_data_i_40));
sg13g2_nand2_2 U140 (.A(data_o_40_), .B(n4321), .Y(n690));
sg13g2_o21ai_1 U141 (.A1(n4328), .A2(n691), .B1(n692), .Y(subbytes_data_i_3));
sg13g2_nand2_2 U142 (.A(data_o_3_), .B(n4321), .Y(n692));
sg13g2_nand3_1 U143 (.A(n1526), .B(n539), .C(n1525), .Y(next_addroundkey_data_reg_29));
sg13g2_nand3_1 U144 (.A(n1521), .B(n540), .C(n1520), .Y(next_addroundkey_data_reg_2));
sg13g2_o21ai_1 U145 (.A1(n4328), .A2(n695), .B1(n696), .Y(subbytes_data_i_38));
sg13g2_nand2_2 U146 (.A(data_o_38_), .B(n4298), .Y(n696));
sg13g2_o21ai_1 U147 (.A1(n4329), .A2(n697), .B1(n698), .Y(subbytes_data_i_37));
sg13g2_nand2_2 U148 (.A(data_o_37_), .B(n4321), .Y(n698));
sg13g2_o21ai_1 U149 (.A1(n4326), .A2(n699), .B1(n700), .Y(subbytes_data_i_36));
sg13g2_nand2_2 U150 (.A(data_o_36_), .B(n4298), .Y(n700));
sg13g2_o21ai_1 U151 (.A1(n4330), .A2(n701), .B1(n702), .Y(subbytes_data_i_35));
sg13g2_nand2_2 U152 (.A(data_o_35_), .B(n4298), .Y(n702));
sg13g2_o21ai_1 U153 (.A1(n4327), .A2(n703), .B1(n704), .Y(subbytes_data_i_34));
sg13g2_nand2_2 U154 (.A(data_o_34_), .B(n4298), .Y(n704));
sg13g2_o21ai_1 U155 (.A1(n4329), .A2(n705), .B1(n706), .Y(subbytes_data_i_33));
sg13g2_nand2_2 U156 (.A(data_o_33_), .B(n4298), .Y(n706));
sg13g2_o21ai_1 U157 (.A1(n4329), .A2(n707), .B1(n708), .Y(subbytes_data_i_32));
sg13g2_nand2_2 U158 (.A(data_o_32_), .B(n4321), .Y(n708));
sg13g2_o21ai_1 U159 (.A1(n4326), .A2(n709), .B1(n710), .Y(subbytes_data_i_31));
sg13g2_nand2_2 U160 (.A(data_o_31_), .B(n4321), .Y(n710));
sg13g2_o21ai_1 U161 (.A1(n4328), .A2(n711), .B1(n712), .Y(subbytes_data_i_30));
sg13g2_nand2_2 U162 (.A(data_o_30_), .B(n4298), .Y(n712));
sg13g2_o21ai_1 U163 (.A1(n4327), .A2(n713), .B1(n714), .Y(subbytes_data_i_2));
sg13g2_nand2_2 U164 (.A(data_o_2_), .B(n4321), .Y(n714));
sg13g2_o21ai_1 U165 (.A1(n4325), .A2(n715), .B1(n716), .Y(subbytes_data_i_29));
sg13g2_nand2_2 U166 (.A(data_o_29_), .B(n4319), .Y(n716));
sg13g2_o21ai_1 U167 (.A1(n4326), .A2(n717), .B1(n718), .Y(subbytes_data_i_28));
sg13g2_nand2_2 U168 (.A(data_o_28_), .B(n4321), .Y(n718));
sg13g2_o21ai_1 U169 (.A1(n4325), .A2(n719), .B1(n720), .Y(subbytes_data_i_27));
sg13g2_nand2_2 U170 (.A(data_o_27_), .B(n4319), .Y(n720));
sg13g2_o21ai_1 U171 (.A1(n4330), .A2(n721), .B1(n722), .Y(subbytes_data_i_26));
sg13g2_nand2_2 U172 (.A(data_o_26_), .B(n4298), .Y(n722));
sg13g2_o21ai_1 U173 (.A1(n4325), .A2(n723), .B1(n724), .Y(subbytes_data_i_25));
sg13g2_nand2_2 U174 (.A(data_o_25_), .B(n4319), .Y(n724));
sg13g2_o21ai_1 U175 (.A1(n4328), .A2(n725), .B1(n726), .Y(subbytes_data_i_24));
sg13g2_nand2_2 U176 (.A(data_o_24_), .B(n4320), .Y(n726));
sg13g2_nand3_1 U177 (.A(n1516), .B(n541), .C(n1515), .Y(next_addroundkey_data_reg_30));
sg13g2_nand2_2 U178 (.A(data_o_23_), .B(n4298), .Y(n728));
sg13g2_o21ai_1 U179 (.A1(n4330), .A2(n729), .B1(n730), .Y(subbytes_data_i_22));
sg13g2_nand2_2 U180 (.A(data_o_22_), .B(n4321), .Y(n730));
sg13g2_o21ai_1 U181 (.A1(n4325), .A2(n731), .B1(n732), .Y(subbytes_data_i_21));
sg13g2_nand2_2 U182 (.A(data_o_21_), .B(n4320), .Y(n732));
sg13g2_o21ai_1 U183 (.A1(n4325), .A2(n733), .B1(n734), .Y(subbytes_data_i_20));
sg13g2_nand2_2 U184 (.A(data_o_20_), .B(n4321), .Y(n734));
sg13g2_o21ai_1 U185 (.A1(n4327), .A2(n735), .B1(n736), .Y(subbytes_data_i_1));
sg13g2_nand2_2 U186 (.A(data_o_1_), .B(n4321), .Y(n736));
sg13g2_o21ai_1 U187 (.A1(n4327), .A2(n737), .B1(n738), .Y(subbytes_data_i_19));
sg13g2_nand2_2 U188 (.A(data_o_19_), .B(n4298), .Y(n738));
sg13g2_o21ai_1 U189 (.A1(n4327), .A2(n739), .B1(n740), .Y(subbytes_data_i_18));
sg13g2_nand2_2 U190 (.A(data_o_18_), .B(n4321), .Y(n740));
sg13g2_o21ai_1 U191 (.A1(n4327), .A2(n741), .B1(n742), .Y(subbytes_data_i_17));
sg13g2_nand2_2 U192 (.A(data_o_17_), .B(n4318), .Y(n742));
sg13g2_o21ai_1 U193 (.A1(n4327), .A2(n743), .B1(n744), .Y(subbytes_data_i_16));
sg13g2_nand2_2 U194 (.A(data_o_16_), .B(n4320), .Y(n744));
sg13g2_nand3_1 U195 (.A(n1511), .B(n542), .C(n1510), .Y(next_addroundkey_data_reg_31));
sg13g2_nand3_1 U196 (.A(n1506), .B(n543), .C(n1505), .Y(next_addroundkey_data_reg_32));
sg13g2_o21ai_1 U197 (.A1(n4327), .A2(n747), .B1(n748), .Y(subbytes_data_i_14));
sg13g2_nand2_2 U198 (.A(data_o_14_), .B(n4298), .Y(n748));
sg13g2_o21ai_1 U199 (.A1(n4327), .A2(n749), .B1(n750), .Y(subbytes_data_i_13));
sg13g2_nand2_2 U200 (.A(data_o_13_), .B(n4321), .Y(n750));
sg13g2_o21ai_1 U201 (.A1(n4327), .A2(n751), .B1(n752), .Y(subbytes_data_i_12));
sg13g2_nand2_2 U202 (.A(data_o_12_), .B(n4321), .Y(n752));
sg13g2_nand3_1 U203 (.A(n1501), .B(n544), .C(n1500), .Y(next_addroundkey_data_reg_33));
sg13g2_nand2_2 U204 (.A(data_o_127_), .B(n4319), .Y(n754));
sg13g2_nand3_1 U205 (.A(n1496), .B(n545), .C(n1495), .Y(next_addroundkey_data_reg_34));
sg13g2_nand2_2 U206 (.A(data_o_126_), .B(n4298), .Y(n756));
sg13g2_o21ai_1 U207 (.A1(n4329), .A2(n757), .B1(n758), .Y(subbytes_data_i_125));
sg13g2_nand2_2 U208 (.A(data_o_125_), .B(n4319), .Y(n758));
sg13g2_nand3_1 U209 (.A(n1491), .B(n546), .C(n1490), .Y(next_addroundkey_data_reg_35));
sg13g2_nand2_2 U210 (.A(data_o_124_), .B(n4298), .Y(n760));
sg13g2_nand3_1 U211 (.A(n1486), .B(n547), .C(n1485), .Y(next_addroundkey_data_reg_36));
sg13g2_nand3_1 U212 (.A(n1481), .B(n548), .C(n1480), .Y(next_addroundkey_data_reg_37));
sg13g2_o21ai_1 U213 (.A1(n4327), .A2(n763), .B1(n764), .Y(subbytes_data_i_122));
sg13g2_nand3_1 U214 (.A(n1476), .B(n556), .C(n1475), .Y(next_addroundkey_data_reg_38));
sg13g2_o21ai_1 U215 (.A1(n4329), .A2(n765), .B1(n766), .Y(subbytes_data_i_121));
sg13g2_nand2_2 U216 (.A(data_o_121_), .B(n4319), .Y(n766));
sg13g2_nand3_1 U217 (.A(n1471), .B(n816), .C(n1470), .Y(next_addroundkey_data_reg_39));
sg13g2_nand2_2 U218 (.A(data_o_120_), .B(n4316), .Y(n768));
sg13g2_o21ai_1 U219 (.A1(n4326), .A2(n769), .B1(n770), .Y(subbytes_data_i_11));
sg13g2_nand2_2 U220 (.A(data_o_11_), .B(n4323), .Y(n770));
sg13g2_o21ai_1 U221 (.A1(n4328), .A2(n771), .B1(n772), .Y(subbytes_data_i_119));
sg13g2_nand2_2 U222 (.A(data_o_119_), .B(n4321), .Y(n772));
sg13g2_o21ai_1 U223 (.A1(n4327), .A2(n773), .B1(n774), .Y(subbytes_data_i_118));
sg13g2_nand3_1 U224 (.A(n1466), .B(n817), .C(n1465), .Y(next_addroundkey_data_reg_3));
sg13g2_o21ai_1 U225 (.A1(n4330), .A2(n775), .B1(n776), .Y(subbytes_data_i_117));
sg13g2_nand2_2 U226 (.A(data_o_117_), .B(n4318), .Y(n776));
sg13g2_o21ai_1 U227 (.A1(n4326), .A2(n777), .B1(n778), .Y(subbytes_data_i_116));
sg13g2_nand2_2 U228 (.A(data_o_116_), .B(n4316), .Y(n778));
sg13g2_o21ai_1 U229 (.A1(n4329), .A2(n779), .B1(n780), .Y(subbytes_data_i_115));
sg13g2_nand2_2 U230 (.A(data_o_115_), .B(n4319), .Y(n780));
sg13g2_o21ai_1 U231 (.A1(n4327), .A2(n781), .B1(n782), .Y(subbytes_data_i_114));
sg13g2_nand2_2 U232 (.A(data_o_114_), .B(n4320), .Y(n782));
sg13g2_o21ai_1 U233 (.A1(n4327), .A2(n783), .B1(n784), .Y(subbytes_data_i_113));
sg13g2_nand2_2 U234 (.A(data_o_113_), .B(n4318), .Y(n784));
sg13g2_o21ai_1 U235 (.A1(n4326), .A2(n785), .B1(n786), .Y(subbytes_data_i_112));
sg13g2_nand2_2 U236 (.A(data_o_112_), .B(n4319), .Y(n786));
sg13g2_nand3_1 U237 (.A(n1461), .B(n819), .C(n1460), .Y(next_addroundkey_data_reg_40));
sg13g2_nand3_1 U238 (.A(n1456), .B(n821), .C(n1455), .Y(next_addroundkey_data_reg_41));
sg13g2_o21ai_1 U239 (.A1(n4325), .A2(n789), .B1(n790), .Y(subbytes_data_i_110));
sg13g2_nand2_2 U240 (.A(data_o_110_), .B(n4317), .Y(n790));
sg13g2_o21ai_1 U241 (.A1(n4326), .A2(n791), .B1(n792), .Y(subbytes_data_i_10));
sg13g2_nand2_2 U242 (.A(data_o_10_), .B(n4317), .Y(n792));
sg13g2_o21ai_1 U243 (.A1(n4329), .A2(n793), .B1(n794), .Y(subbytes_data_i_109));
sg13g2_nand2_2 U244 (.A(data_o_109_), .B(n4317), .Y(n794));
sg13g2_o21ai_1 U245 (.A1(n4326), .A2(n795), .B1(n796), .Y(subbytes_data_i_108));
sg13g2_nand2_2 U246 (.A(data_o_108_), .B(n4319), .Y(n796));
sg13g2_o21ai_1 U247 (.A1(n4325), .A2(n797), .B1(n798), .Y(subbytes_data_i_107));
sg13g2_nand2_2 U248 (.A(data_o_107_), .B(n4319), .Y(n798));
sg13g2_o21ai_1 U249 (.A1(n4326), .A2(n799), .B1(n800), .Y(subbytes_data_i_106));
sg13g2_nand2_2 U250 (.A(data_o_106_), .B(n4321), .Y(n800));
sg13g2_o21ai_1 U251 (.A1(n4326), .A2(n801), .B1(n802), .Y(subbytes_data_i_105));
sg13g2_nand2_2 U252 (.A(data_o_105_), .B(n4321), .Y(n802));
sg13g2_o21ai_1 U253 (.A1(n4325), .A2(n803), .B1(n804), .Y(subbytes_data_i_104));
sg13g2_nand2_2 U254 (.A(data_o_104_), .B(n4318), .Y(n804));
sg13g2_o21ai_1 U255 (.A1(n4330), .A2(n805), .B1(n806), .Y(subbytes_data_i_103));
sg13g2_nand2_2 U256 (.A(data_o_103_), .B(n4316), .Y(n806));
sg13g2_o21ai_1 U257 (.A1(n4330), .A2(n807), .B1(n808), .Y(subbytes_data_i_102));
sg13g2_nand2_2 U258 (.A(data_o_102_), .B(n4320), .Y(n808));
sg13g2_o21ai_1 U259 (.A1(n4328), .A2(n809), .B1(n810), .Y(subbytes_data_i_101));
sg13g2_nand2_2 U260 (.A(data_o_101_), .B(n4319), .Y(n810));
sg13g2_o21ai_1 U261 (.A1(n4328), .A2(n811), .B1(n812), .Y(subbytes_data_i_100));
sg13g2_nand2_2 U262 (.A(data_o_100_), .B(n4316), .Y(n812));
sg13g2_o21ai_1 U263 (.A1(n4326), .A2(n813), .B1(n814), .Y(subbytes_data_i_0));
sg13g2_nand2_2 U264 (.A(data_o_0_), .B(n4321), .Y(n814));
sg13g2_nand3_1 U265 (.A(n1451), .B(n823), .C(n1450), .Y(next_addroundkey_data_reg_42));
sg13g2_nand3_1 U266 (.A(n1446), .B(n825), .C(n1445), .Y(next_addroundkey_data_reg_43));
sg13g2_inv_4 U267 (.A(subbytes_sbox_decrypt_o), .Y(n815));
sg13g2_nand3_1 U268 (.A(n1441), .B(n827), .C(n1440), .Y(next_addroundkey_data_reg_44));
sg13g2_nand3_1 U269 (.A(n1436), .B(n829), .C(n1435), .Y(next_addroundkey_data_reg_45));
sg13g2_nand3_1 U270 (.A(n1431), .B(n831), .C(n1430), .Y(next_addroundkey_data_reg_46));
sg13g2_nand3_1 U271 (.A(n1426), .B(n833), .C(n1425), .Y(next_addroundkey_data_reg_47));
sg13g2_nand3_1 U272 (.A(n1421), .B(n842), .C(n1420), .Y(next_addroundkey_data_reg_48));
sg13g2_nand3_1 U273 (.A(n1416), .B(n854), .C(n1415), .Y(next_addroundkey_data_reg_49));
sg13g2_nand3_1 U274 (.A(n1411), .B(n1110), .C(n1410), .Y(next_addroundkey_data_reg_4));
sg13g2_nand3_1 U275 (.A(n1406), .B(n1111), .C(n1405), .Y(next_addroundkey_data_reg_50));
sg13g2_nand3_1 U276 (.A(n1401), .B(n1112), .C(n1400), .Y(next_addroundkey_data_reg_51));
sg13g2_nand3_1 U277 (.A(n1396), .B(n1113), .C(n1395), .Y(next_addroundkey_data_reg_52));
sg13g2_nand3_1 U278 (.A(n1391), .B(n1114), .C(n1390), .Y(next_addroundkey_data_reg_53));
sg13g2_nand3_1 U279 (.A(n1386), .B(n1125), .C(n1385), .Y(next_addroundkey_data_reg_54));
sg13g2_nand3_1 U280 (.A(n1381), .B(n1130), .C(n1380), .Y(next_addroundkey_data_reg_55));
sg13g2_nand3_1 U281 (.A(n1376), .B(n1137), .C(n1375), .Y(next_addroundkey_data_reg_56));
sg13g2_nand3_1 U282 (.A(n1371), .B(n1138), .C(n1370), .Y(next_addroundkey_data_reg_57));
sg13g2_nand3_1 U283 (.A(n1366), .B(n1906), .C(n1365), .Y(next_addroundkey_data_reg_58));
sg13g2_nand3_1 U284 (.A(n1361), .B(n1908), .C(n1360), .Y(next_addroundkey_data_reg_59));
sg13g2_nand3_1 U285 (.A(n1356), .B(n1915), .C(n1355), .Y(next_addroundkey_data_reg_5));
sg13g2_nand3_1 U286 (.A(n1351), .B(n1916), .C(n1350), .Y(next_addroundkey_data_reg_60));
sg13g2_nand3_1 U287 (.A(n1346), .B(n2173), .C(n1345), .Y(next_addroundkey_data_reg_61));
sg13g2_nand3_1 U288 (.A(n1341), .B(n2236), .C(n1340), .Y(next_addroundkey_data_reg_62));
sg13g2_nand3_1 U289 (.A(n1336), .B(n2237), .C(n1335), .Y(next_addroundkey_data_reg_63));
sg13g2_nand3_1 U290 (.A(n1331), .B(n2238), .C(n1330), .Y(next_addroundkey_data_reg_64));
sg13g2_nand3_1 U291 (.A(n1326), .B(n2239), .C(n1325), .Y(next_addroundkey_data_reg_65));
sg13g2_nand3_1 U292 (.A(n1321), .B(n2240), .C(n1320), .Y(next_addroundkey_data_reg_66));
sg13g2_nand2_2 U293 (.A(n835), .B(n836), .Y(n834));
sg13g2_o21ai_1 U294 (.A1(n837), .A2(N1), .B1(n838), .Y(n836));
sg13g2_nand2_2 U295 (.A(N175), .B(n837), .Y(n838));
sg13g2_nand3_1 U296 (.A(n1316), .B(n3524), .C(n1315), .Y(next_addroundkey_data_reg_67));
sg13g2_nand2_2 U297 (.A(n835), .B(n840), .Y(n839));
sg13g2_o21ai_1 U298 (.A1(net47628), .A2(n837), .B1(n841), .Y(n840));
sg13g2_nand2_2 U299 (.A(N174), .B(n837), .Y(n841));
sg13g2_nand2_2 U300 (.A(n4315), .B(n843), .Y(n837));
sg13g2_nand3_1 U301 (.A(n1311), .B(n3658), .C(n1310), .Y(next_addroundkey_data_reg_68));
sg13g2_a21oi_2 U302 (.A1(n844), .A2(n845), .B1(n846), .Y(next_round_1));
sg13g2_nand3_1 U303 (.A(n1306), .B(n3659), .C(n1305), .Y(next_addroundkey_data_reg_69));
sg13g2_nand2_2 U304 (.A(three_1), .B(n848), .Y(n844));
sg13g2_inv_4 U305 (.A(n847), .Y(n848));
sg13g2_nor2_2 U306 (.A(n846), .B(n849), .Y(next_round_0));
sg13g2_xnor2_1 U307 (.A(three_0), .B(n847), .Y(n849));
sg13g2_nor2_2 U308 (.A(n850), .B(n851), .Y(n847));
sg13g2_o21ai_1 U309 (.A1(net24693), .A2(n852), .B1(n853), .Y(next_last_key_half_9));
sg13g2_a21oi_2 U310 (.A1(last_key_half_9), .A2(net26864), .B1(n855), .Y(n853));
sg13g2_inv_4 U311 (.A(n856), .Y(n855));
sg13g2_nand2_2 U312 (.A(n857), .B(keysched_new_key_o_9), .Y(n856));
sg13g2_o21ai_1 U313 (.A1(net24693), .A2(n858), .B1(n859), .Y(next_last_key_half_8));
sg13g2_a21oi_2 U314 (.A1(last_key_half_8), .A2(net26864), .B1(n860), .Y(n859));
sg13g2_inv_4 U315 (.A(n861), .Y(n860));
sg13g2_nand2_2 U316 (.A(n857), .B(keysched_new_key_o_8), .Y(n861));
sg13g2_o21ai_1 U317 (.A1(net24693), .A2(n862), .B1(n863), .Y(next_last_key_half_7));
sg13g2_a21oi_2 U318 (.A1(last_key_half_7), .A2(net26864), .B1(n864), .Y(n863));
sg13g2_inv_4 U319 (.A(n865), .Y(n864));
sg13g2_nand2_2 U320 (.A(n857), .B(keysched_new_key_o_7), .Y(n865));
sg13g2_o21ai_1 U321 (.A1(net24693), .A2(n866), .B1(n867), .Y(next_last_key_half_6));
sg13g2_a21oi_2 U322 (.A1(last_key_half_6), .A2(net26864), .B1(n868), .Y(n867));
sg13g2_inv_4 U323 (.A(n869), .Y(n868));
sg13g2_nand2_2 U324 (.A(n857), .B(keysched_new_key_o_6), .Y(n869));
sg13g2_o21ai_1 U325 (.A1(net24693), .A2(n870), .B1(n871), .Y(next_last_key_half_63));
sg13g2_a21oi_2 U326 (.A1(last_key_half_63), .A2(net26864), .B1(n872), .Y(n871));
sg13g2_inv_4 U327 (.A(n873), .Y(n872));
sg13g2_nand2_2 U328 (.A(n857), .B(keysched_new_key_o_63), .Y(n873));
sg13g2_o21ai_1 U329 (.A1(net24693), .A2(n874), .B1(n875), .Y(next_last_key_half_62));
sg13g2_a21oi_2 U330 (.A1(last_key_half_62), .A2(net26864), .B1(n876), .Y(n875));
sg13g2_inv_4 U331 (.A(n877), .Y(n876));
sg13g2_nand2_2 U332 (.A(n857), .B(keysched_new_key_o_62), .Y(n877));
sg13g2_o21ai_1 U333 (.A1(net24693), .A2(n878), .B1(n879), .Y(next_last_key_half_61));
sg13g2_a21oi_2 U334 (.A1(last_key_half_61), .A2(net26864), .B1(n880), .Y(n879));
sg13g2_inv_4 U335 (.A(n881), .Y(n880));
sg13g2_nand2_2 U336 (.A(n857), .B(keysched_new_key_o_61), .Y(n881));
sg13g2_o21ai_1 U337 (.A1(net24693), .A2(n882), .B1(n883), .Y(next_last_key_half_60));
sg13g2_a21oi_2 U338 (.A1(last_key_half_60), .A2(net26864), .B1(n884), .Y(n883));
sg13g2_inv_4 U339 (.A(n885), .Y(n884));
sg13g2_nand2_2 U340 (.A(n857), .B(keysched_new_key_o_60), .Y(n885));
sg13g2_o21ai_1 U341 (.A1(net24693), .A2(n886), .B1(n887), .Y(next_last_key_half_5));
sg13g2_a21oi_2 U342 (.A1(last_key_half_5), .A2(net26864), .B1(n888), .Y(n887));
sg13g2_inv_4 U343 (.A(n889), .Y(n888));
sg13g2_nand2_2 U344 (.A(n857), .B(keysched_new_key_o_5), .Y(n889));
sg13g2_o21ai_1 U345 (.A1(net24693), .A2(n890), .B1(n891), .Y(next_last_key_half_59));
sg13g2_a21oi_2 U346 (.A1(last_key_half_59), .A2(net26864), .B1(n892), .Y(n891));
sg13g2_inv_4 U347 (.A(n893), .Y(n892));
sg13g2_nand2_2 U348 (.A(n857), .B(keysched_new_key_o_59), .Y(n893));
sg13g2_o21ai_1 U349 (.A1(net24693), .A2(n894), .B1(n895), .Y(next_last_key_half_58));
sg13g2_a21oi_2 U350 (.A1(last_key_half_58), .A2(net26864), .B1(n896), .Y(n895));
sg13g2_inv_4 U351 (.A(n897), .Y(n896));
sg13g2_nand2_2 U352 (.A(n857), .B(keysched_new_key_o_58), .Y(n897));
sg13g2_o21ai_1 U353 (.A1(net24693), .A2(n898), .B1(n899), .Y(next_last_key_half_57));
sg13g2_a21oi_2 U354 (.A1(last_key_half_57), .A2(net26864), .B1(n900), .Y(n899));
sg13g2_inv_4 U355 (.A(n901), .Y(n900));
sg13g2_nand2_2 U356 (.A(n857), .B(keysched_new_key_o_57), .Y(n901));
sg13g2_o21ai_1 U357 (.A1(net24693), .A2(n902), .B1(n903), .Y(next_last_key_half_56));
sg13g2_a21oi_2 U358 (.A1(last_key_half_56), .A2(net26864), .B1(n904), .Y(n903));
sg13g2_inv_4 U359 (.A(n905), .Y(n904));
sg13g2_nand2_2 U360 (.A(n857), .B(keysched_new_key_o_56), .Y(n905));
sg13g2_o21ai_1 U361 (.A1(net24693), .A2(n906), .B1(n907), .Y(next_last_key_half_55));
sg13g2_a21oi_2 U362 (.A1(last_key_half_55), .A2(net26864), .B1(n908), .Y(n907));
sg13g2_inv_4 U363 (.A(n909), .Y(n908));
sg13g2_nand2_2 U364 (.A(n857), .B(keysched_new_key_o_55), .Y(n909));
sg13g2_o21ai_1 U365 (.A1(net24693), .A2(n910), .B1(n911), .Y(next_last_key_half_54));
sg13g2_a21oi_2 U366 (.A1(last_key_half_54), .A2(net26864), .B1(n912), .Y(n911));
sg13g2_inv_4 U367 (.A(n913), .Y(n912));
sg13g2_nand2_2 U368 (.A(n857), .B(keysched_new_key_o_54), .Y(n913));
sg13g2_o21ai_1 U369 (.A1(net24693), .A2(n914), .B1(n915), .Y(next_last_key_half_53));
sg13g2_a21oi_2 U370 (.A1(last_key_half_53), .A2(net26864), .B1(n916), .Y(n915));
sg13g2_inv_4 U371 (.A(n917), .Y(n916));
sg13g2_nand2_2 U372 (.A(n857), .B(keysched_new_key_o_53), .Y(n917));
sg13g2_o21ai_1 U373 (.A1(net24693), .A2(n918), .B1(n919), .Y(next_last_key_half_52));
sg13g2_a21oi_2 U374 (.A1(last_key_half_52), .A2(net26864), .B1(n920), .Y(n919));
sg13g2_inv_4 U375 (.A(n921), .Y(n920));
sg13g2_nand2_2 U376 (.A(n857), .B(keysched_new_key_o_52), .Y(n921));
sg13g2_o21ai_1 U377 (.A1(net24693), .A2(n922), .B1(n923), .Y(next_last_key_half_51));
sg13g2_a21oi_2 U378 (.A1(last_key_half_51), .A2(net26864), .B1(n924), .Y(n923));
sg13g2_inv_4 U379 (.A(n925), .Y(n924));
sg13g2_nand2_2 U380 (.A(n857), .B(keysched_new_key_o_51), .Y(n925));
sg13g2_o21ai_1 U381 (.A1(net24693), .A2(n926), .B1(n927), .Y(next_last_key_half_50));
sg13g2_a21oi_2 U382 (.A1(last_key_half_50), .A2(net26864), .B1(n928), .Y(n927));
sg13g2_inv_4 U383 (.A(n929), .Y(n928));
sg13g2_nand2_2 U384 (.A(n857), .B(keysched_new_key_o_50), .Y(n929));
sg13g2_o21ai_1 U385 (.A1(net24693), .A2(n930), .B1(n931), .Y(next_last_key_half_4));
sg13g2_a21oi_2 U386 (.A1(last_key_half_4), .A2(net26864), .B1(n932), .Y(n931));
sg13g2_inv_4 U387 (.A(n933), .Y(n932));
sg13g2_nand2_2 U388 (.A(n857), .B(keysched_new_key_o_4), .Y(n933));
sg13g2_o21ai_1 U389 (.A1(net24693), .A2(n934), .B1(n935), .Y(next_last_key_half_49));
sg13g2_a21oi_2 U390 (.A1(last_key_half_49), .A2(net26864), .B1(n936), .Y(n935));
sg13g2_inv_4 U391 (.A(n937), .Y(n936));
sg13g2_nand2_2 U392 (.A(n857), .B(keysched_new_key_o_49), .Y(n937));
sg13g2_nand3_1 U393 (.A(n1301), .B(n3660), .C(n1300), .Y(next_addroundkey_data_reg_6));
sg13g2_a21oi_2 U394 (.A1(last_key_half_48), .A2(net26864), .B1(n940), .Y(n939));
sg13g2_inv_4 U395 (.A(n941), .Y(n940));
sg13g2_nand2_2 U396 (.A(n857), .B(keysched_new_key_o_48), .Y(n941));
sg13g2_o21ai_1 U397 (.A1(net24693), .A2(n942), .B1(n943), .Y(next_last_key_half_47));
sg13g2_a21oi_2 U398 (.A1(last_key_half_47), .A2(net26864), .B1(n944), .Y(n943));
sg13g2_inv_4 U399 (.A(n945), .Y(n944));
sg13g2_nand2_2 U400 (.A(n857), .B(keysched_new_key_o_47), .Y(n945));
sg13g2_nand3_1 U401 (.A(n1296), .B(n3661), .C(n1295), .Y(next_addroundkey_data_reg_70));
sg13g2_nand3_1 U402 (.A(n1291), .B(n3662), .C(n1290), .Y(next_addroundkey_data_reg_71));
sg13g2_inv_4 U403 (.A(n949), .Y(n948));
sg13g2_nand2_2 U404 (.A(n857), .B(keysched_new_key_o_46), .Y(n949));
sg13g2_o21ai_1 U405 (.A1(net24693), .A2(n950), .B1(n951), .Y(next_last_key_half_45));
sg13g2_a21oi_2 U406 (.A1(last_key_half_45), .A2(net26864), .B1(n952), .Y(n951));
sg13g2_inv_4 U407 (.A(n953), .Y(n952));
sg13g2_nand2_2 U408 (.A(n857), .B(keysched_new_key_o_45), .Y(n953));
sg13g2_o21ai_1 U409 (.A1(net24693), .A2(n954), .B1(n955), .Y(next_last_key_half_44));
sg13g2_a21oi_2 U410 (.A1(last_key_half_44), .A2(net26864), .B1(n956), .Y(n955));
sg13g2_inv_4 U411 (.A(n957), .Y(n956));
sg13g2_nand2_2 U412 (.A(n857), .B(keysched_new_key_o_44), .Y(n957));
sg13g2_o21ai_1 U413 (.A1(net24693), .A2(n958), .B1(n959), .Y(next_last_key_half_43));
sg13g2_a21oi_2 U414 (.A1(last_key_half_43), .A2(net26864), .B1(n960), .Y(n959));
sg13g2_inv_4 U415 (.A(n961), .Y(n960));
sg13g2_nand2_2 U416 (.A(n857), .B(keysched_new_key_o_43), .Y(n961));
sg13g2_o21ai_1 U417 (.A1(net24693), .A2(n962), .B1(n963), .Y(next_last_key_half_42));
sg13g2_a21oi_2 U418 (.A1(last_key_half_42), .A2(net26864), .B1(n964), .Y(n963));
sg13g2_inv_4 U419 (.A(n965), .Y(n964));
sg13g2_nand2_2 U420 (.A(n857), .B(keysched_new_key_o_42), .Y(n965));
sg13g2_o21ai_1 U421 (.A1(net24693), .A2(n966), .B1(n967), .Y(next_last_key_half_41));
sg13g2_a21oi_2 U422 (.A1(last_key_half_41), .A2(net26864), .B1(n968), .Y(n967));
sg13g2_inv_4 U423 (.A(n969), .Y(n968));
sg13g2_nand2_2 U424 (.A(n857), .B(keysched_new_key_o_41), .Y(n969));
sg13g2_o21ai_1 U425 (.A1(net24693), .A2(n970), .B1(n971), .Y(next_last_key_half_40));
sg13g2_a21oi_2 U426 (.A1(last_key_half_40), .A2(net26864), .B1(n972), .Y(n971));
sg13g2_inv_4 U427 (.A(n973), .Y(n972));
sg13g2_nand2_2 U428 (.A(n857), .B(keysched_new_key_o_40), .Y(n973));
sg13g2_o21ai_1 U429 (.A1(net24693), .A2(n974), .B1(n975), .Y(next_last_key_half_3));
sg13g2_a21oi_2 U430 (.A1(last_key_half_3), .A2(net26864), .B1(n976), .Y(n975));
sg13g2_inv_4 U431 (.A(n977), .Y(n976));
sg13g2_nand2_2 U432 (.A(n857), .B(keysched_new_key_o_3), .Y(n977));
sg13g2_o21ai_1 U433 (.A1(net24693), .A2(n978), .B1(n979), .Y(next_last_key_half_39));
sg13g2_a21oi_2 U434 (.A1(last_key_half_39), .A2(net26864), .B1(n980), .Y(n979));
sg13g2_inv_4 U435 (.A(n981), .Y(n980));
sg13g2_nand2_2 U436 (.A(n857), .B(keysched_new_key_o_39), .Y(n981));
sg13g2_o21ai_1 U437 (.A1(net24693), .A2(n982), .B1(n983), .Y(next_last_key_half_38));
sg13g2_a21oi_2 U438 (.A1(last_key_half_38), .A2(net26864), .B1(n984), .Y(n983));
sg13g2_inv_4 U439 (.A(n985), .Y(n984));
sg13g2_nand2_2 U440 (.A(n857), .B(keysched_new_key_o_38), .Y(n985));
sg13g2_o21ai_1 U441 (.A1(net24693), .A2(n986), .B1(n987), .Y(next_last_key_half_37));
sg13g2_a21oi_2 U442 (.A1(last_key_half_37), .A2(net26864), .B1(n988), .Y(n987));
sg13g2_inv_4 U443 (.A(n989), .Y(n988));
sg13g2_nand2_2 U444 (.A(n857), .B(keysched_new_key_o_37), .Y(n989));
sg13g2_o21ai_1 U445 (.A1(net24693), .A2(n990), .B1(n991), .Y(next_last_key_half_36));
sg13g2_a21oi_2 U446 (.A1(last_key_half_36), .A2(net26864), .B1(n992), .Y(n991));
sg13g2_inv_4 U447 (.A(n993), .Y(n992));
sg13g2_nand2_2 U448 (.A(n857), .B(keysched_new_key_o_36), .Y(n993));
sg13g2_o21ai_1 U449 (.A1(net24693), .A2(n994), .B1(n995), .Y(next_last_key_half_35));
sg13g2_a21oi_2 U450 (.A1(last_key_half_35), .A2(net26864), .B1(n996), .Y(n995));
sg13g2_inv_4 U451 (.A(n997), .Y(n996));
sg13g2_nand2_2 U452 (.A(n857), .B(keysched_new_key_o_35), .Y(n997));
sg13g2_o21ai_1 U453 (.A1(net24693), .A2(n998), .B1(n999), .Y(next_last_key_half_34));
sg13g2_a21oi_2 U454 (.A1(last_key_half_34), .A2(net26864), .B1(n1000), .Y(n999));
sg13g2_inv_4 U455 (.A(n1001), .Y(n1000));
sg13g2_nand2_2 U456 (.A(n857), .B(keysched_new_key_o_34), .Y(n1001));
sg13g2_o21ai_1 U457 (.A1(net24693), .A2(n1002), .B1(n1003), .Y(next_last_key_half_33));
sg13g2_a21oi_2 U458 (.A1(last_key_half_33), .A2(net26864), .B1(n1004), .Y(n1003));
sg13g2_inv_4 U459 (.A(n1005), .Y(n1004));
sg13g2_nand2_2 U460 (.A(n857), .B(keysched_new_key_o_33), .Y(n1005));
sg13g2_o21ai_1 U461 (.A1(net24693), .A2(n1006), .B1(n1007), .Y(next_last_key_half_32));
sg13g2_a21oi_2 U462 (.A1(last_key_half_32), .A2(net26864), .B1(n1008), .Y(n1007));
sg13g2_inv_4 U463 (.A(n1009), .Y(n1008));
sg13g2_nand2_2 U464 (.A(n857), .B(keysched_new_key_o_32), .Y(n1009));
sg13g2_o21ai_1 U465 (.A1(net24693), .A2(n1010), .B1(n1011), .Y(next_last_key_half_31));
sg13g2_a21oi_2 U466 (.A1(last_key_half_31), .A2(net26864), .B1(n1012), .Y(n1011));
sg13g2_inv_4 U467 (.A(n1013), .Y(n1012));
sg13g2_nand2_2 U468 (.A(n857), .B(keysched_new_key_o_31), .Y(n1013));
sg13g2_o21ai_1 U469 (.A1(net24693), .A2(n1014), .B1(n1015), .Y(next_last_key_half_30));
sg13g2_a21oi_2 U470 (.A1(last_key_half_30), .A2(net26864), .B1(n1016), .Y(n1015));
sg13g2_inv_4 U471 (.A(n1017), .Y(n1016));
sg13g2_nand2_2 U472 (.A(n857), .B(keysched_new_key_o_30), .Y(n1017));
sg13g2_o21ai_1 U473 (.A1(net24693), .A2(n1018), .B1(n1019), .Y(next_last_key_half_2));
sg13g2_a21oi_2 U474 (.A1(last_key_half_2), .A2(net26864), .B1(n1020), .Y(n1019));
sg13g2_inv_4 U475 (.A(n1021), .Y(n1020));
sg13g2_nand2_2 U476 (.A(n857), .B(keysched_new_key_o_2), .Y(n1021));
sg13g2_o21ai_1 U477 (.A1(net24693), .A2(n1022), .B1(n1023), .Y(next_last_key_half_29));
sg13g2_a21oi_2 U478 (.A1(last_key_half_29), .A2(net26864), .B1(n1024), .Y(n1023));
sg13g2_inv_4 U479 (.A(n1025), .Y(n1024));
sg13g2_nand2_2 U480 (.A(n857), .B(keysched_new_key_o_29), .Y(n1025));
sg13g2_o21ai_1 U481 (.A1(net24693), .A2(n1026), .B1(n1027), .Y(next_last_key_half_28));
sg13g2_a21oi_2 U482 (.A1(last_key_half_28), .A2(net26864), .B1(n1028), .Y(n1027));
sg13g2_inv_4 U483 (.A(n1029), .Y(n1028));
sg13g2_nand2_2 U484 (.A(n857), .B(keysched_new_key_o_28), .Y(n1029));
sg13g2_o21ai_1 U485 (.A1(net24693), .A2(n1030), .B1(n1031), .Y(next_last_key_half_27));
sg13g2_a21oi_2 U486 (.A1(last_key_half_27), .A2(net26864), .B1(n1032), .Y(n1031));
sg13g2_inv_4 U487 (.A(n1033), .Y(n1032));
sg13g2_nand2_2 U488 (.A(n857), .B(keysched_new_key_o_27), .Y(n1033));
sg13g2_o21ai_1 U489 (.A1(net24693), .A2(n1034), .B1(n1035), .Y(next_last_key_half_26));
sg13g2_a21oi_2 U490 (.A1(last_key_half_26), .A2(net26864), .B1(n1036), .Y(n1035));
sg13g2_inv_4 U491 (.A(n1037), .Y(n1036));
sg13g2_nand2_2 U492 (.A(n857), .B(keysched_new_key_o_26), .Y(n1037));
sg13g2_o21ai_1 U493 (.A1(net24693), .A2(n1038), .B1(n1039), .Y(next_last_key_half_25));
sg13g2_a21oi_2 U494 (.A1(last_key_half_25), .A2(net26864), .B1(n1040), .Y(n1039));
sg13g2_inv_4 U495 (.A(n1041), .Y(n1040));
sg13g2_nand2_2 U496 (.A(n857), .B(keysched_new_key_o_25), .Y(n1041));
sg13g2_o21ai_1 U497 (.A1(net24693), .A2(n1042), .B1(n1043), .Y(next_last_key_half_24));
sg13g2_a21oi_2 U498 (.A1(last_key_half_24), .A2(net26864), .B1(n1044), .Y(n1043));
sg13g2_inv_4 U499 (.A(n1045), .Y(n1044));
sg13g2_nand2_2 U500 (.A(n857), .B(keysched_new_key_o_24), .Y(n1045));
sg13g2_o21ai_1 U501 (.A1(net24693), .A2(n1046), .B1(n1047), .Y(next_last_key_half_23));
sg13g2_a21oi_2 U502 (.A1(last_key_half_23), .A2(net26864), .B1(n1048), .Y(n1047));
sg13g2_inv_4 U503 (.A(n1049), .Y(n1048));
sg13g2_nand2_2 U504 (.A(n857), .B(keysched_new_key_o_23), .Y(n1049));
sg13g2_o21ai_1 U505 (.A1(net24693), .A2(n1050), .B1(n1051), .Y(next_last_key_half_22));
sg13g2_a21oi_2 U506 (.A1(last_key_half_22), .A2(net26864), .B1(n1052), .Y(n1051));
sg13g2_inv_4 U507 (.A(n1053), .Y(n1052));
sg13g2_nand2_2 U508 (.A(n857), .B(keysched_new_key_o_22), .Y(n1053));
sg13g2_o21ai_1 U509 (.A1(net24693), .A2(n1054), .B1(n1055), .Y(next_last_key_half_21));
sg13g2_a21oi_2 U510 (.A1(last_key_half_21), .A2(net26864), .B1(n1056), .Y(n1055));
sg13g2_inv_4 U511 (.A(n1057), .Y(n1056));
sg13g2_nand2_2 U512 (.A(n857), .B(keysched_new_key_o_21), .Y(n1057));
sg13g2_o21ai_1 U513 (.A1(net24693), .A2(n1058), .B1(n1059), .Y(next_last_key_half_20));
sg13g2_a21oi_2 U514 (.A1(last_key_half_20), .A2(net26864), .B1(n1060), .Y(n1059));
sg13g2_inv_4 U515 (.A(n1061), .Y(n1060));
sg13g2_nand2_2 U516 (.A(n857), .B(keysched_new_key_o_20), .Y(n1061));
sg13g2_o21ai_1 U517 (.A1(net24693), .A2(n1062), .B1(n1063), .Y(next_last_key_half_1));
sg13g2_a21oi_2 U518 (.A1(last_key_half_1), .A2(net26864), .B1(n1064), .Y(n1063));
sg13g2_inv_4 U519 (.A(n1065), .Y(n1064));
sg13g2_nand2_2 U520 (.A(n857), .B(keysched_new_key_o_1), .Y(n1065));
sg13g2_o21ai_1 U521 (.A1(net24693), .A2(n1066), .B1(n1067), .Y(next_last_key_half_19));
sg13g2_a21oi_2 U522 (.A1(last_key_half_19), .A2(net26864), .B1(n1068), .Y(n1067));
sg13g2_inv_4 U523 (.A(n1069), .Y(n1068));
sg13g2_nand2_2 U524 (.A(n857), .B(keysched_new_key_o_19), .Y(n1069));
sg13g2_o21ai_1 U525 (.A1(net24693), .A2(n1070), .B1(n1071), .Y(next_last_key_half_18));
sg13g2_a21oi_2 U526 (.A1(last_key_half_18), .A2(net26864), .B1(n1072), .Y(n1071));
sg13g2_inv_4 U527 (.A(n1073), .Y(n1072));
sg13g2_nand2_2 U528 (.A(n857), .B(keysched_new_key_o_18), .Y(n1073));
sg13g2_o21ai_1 U529 (.A1(net24693), .A2(n1074), .B1(n1075), .Y(next_last_key_half_17));
sg13g2_a21oi_2 U530 (.A1(last_key_half_17), .A2(net26864), .B1(n1076), .Y(n1075));
sg13g2_inv_4 U531 (.A(n1077), .Y(n1076));
sg13g2_nand2_2 U532 (.A(n857), .B(keysched_new_key_o_17), .Y(n1077));
sg13g2_o21ai_1 U533 (.A1(net24693), .A2(n1078), .B1(n1079), .Y(next_last_key_half_16));
sg13g2_a21oi_2 U534 (.A1(last_key_half_16), .A2(net26864), .B1(n1080), .Y(n1079));
sg13g2_inv_4 U535 (.A(n1081), .Y(n1080));
sg13g2_nand2_2 U536 (.A(n857), .B(keysched_new_key_o_16), .Y(n1081));
sg13g2_o21ai_1 U537 (.A1(net24693), .A2(n1082), .B1(n1083), .Y(next_last_key_half_15));
sg13g2_a21oi_2 U538 (.A1(last_key_half_15), .A2(net26864), .B1(n1084), .Y(n1083));
sg13g2_inv_4 U539 (.A(n1085), .Y(n1084));
sg13g2_nand2_2 U540 (.A(n857), .B(keysched_new_key_o_15), .Y(n1085));
sg13g2_o21ai_1 U541 (.A1(net24693), .A2(n1086), .B1(n1087), .Y(next_last_key_half_14));
sg13g2_a21oi_2 U542 (.A1(last_key_half_14), .A2(net26864), .B1(n1088), .Y(n1087));
sg13g2_inv_4 U543 (.A(n1089), .Y(n1088));
sg13g2_nand2_2 U544 (.A(n857), .B(keysched_new_key_o_14), .Y(n1089));
sg13g2_o21ai_1 U545 (.A1(net24693), .A2(n1090), .B1(n1091), .Y(next_last_key_half_13));
sg13g2_a21oi_2 U546 (.A1(last_key_half_13), .A2(net26864), .B1(n1092), .Y(n1091));
sg13g2_inv_4 U547 (.A(n1093), .Y(n1092));
sg13g2_nand2_2 U548 (.A(n857), .B(keysched_new_key_o_13), .Y(n1093));
sg13g2_o21ai_1 U549 (.A1(net24693), .A2(n1094), .B1(n1095), .Y(next_last_key_half_12));
sg13g2_a21oi_2 U550 (.A1(last_key_half_12), .A2(net26864), .B1(n1096), .Y(n1095));
sg13g2_inv_4 U551 (.A(n1097), .Y(n1096));
sg13g2_nand2_2 U552 (.A(n857), .B(keysched_new_key_o_12), .Y(n1097));
sg13g2_o21ai_1 U553 (.A1(net24693), .A2(n1098), .B1(n1099), .Y(next_last_key_half_11));
sg13g2_a21oi_2 U554 (.A1(last_key_half_11), .A2(net26864), .B1(n1100), .Y(n1099));
sg13g2_inv_4 U555 (.A(n1101), .Y(n1100));
sg13g2_nand2_2 U556 (.A(n857), .B(keysched_new_key_o_11), .Y(n1101));
sg13g2_o21ai_1 U557 (.A1(net24693), .A2(n1102), .B1(n1103), .Y(next_last_key_half_10));
sg13g2_a21oi_2 U558 (.A1(last_key_half_10), .A2(net26864), .B1(n1104), .Y(n1103));
sg13g2_inv_4 U559 (.A(n1105), .Y(n1104));
sg13g2_nand2_2 U560 (.A(n857), .B(keysched_new_key_o_10), .Y(n1105));
sg13g2_o21ai_1 U561 (.A1(net24693), .A2(n1106), .B1(n1107), .Y(next_last_key_half_0));
sg13g2_a21oi_2 U562 (.A1(last_key_half_0), .A2(net26864), .B1(n1108), .Y(n1107));
sg13g2_inv_4 U563 (.A(n1109), .Y(n1108));
sg13g2_nand2_2 U564 (.A(n857), .B(keysched_new_key_o_0), .Y(n1109));
sg13g2_nand3_1 U565 (.A(n1286), .B(n3663), .C(n1285), .Y(next_addroundkey_data_reg_72));
sg13g2_nand3_1 U566 (.A(n1281), .B(n3664), .C(n1280), .Y(next_addroundkey_data_reg_73));
sg13g2_nand3_1 U567 (.A(n1276), .B(n3665), .C(n1275), .Y(next_addroundkey_data_reg_74));
sg13g2_o21ai_1 U568 (.A1(n1117), .A2(n850), .B1(n835), .Y(n1116));
sg13g2_inv_4 U569 (.A(n846), .Y(n835));
sg13g2_nand2_2 U570 (.A(state), .B(n1118), .Y(n846));
sg13g2_inv_4 U571 (.A(n843), .Y(n850));
sg13g2_a21oi_2 U572 (.A1(n4315), .A2(n1115), .B1(N313), .Y(n1117));
sg13g2_nand3_1 U573 (.A(n1271), .B(n3666), .C(n1270), .Y(next_addroundkey_data_reg_75));
sg13g2_inv_4 U574 (.A(n1119), .Y(next_addroundkey_round_3));
sg13g2_a21oi_2 U575 (.A1(n1120), .A2(N1538), .B1(n1121), .Y(n1119));
sg13g2_nand3_1 U576 (.A(n1266), .B(n3667), .C(n1265), .Y(next_addroundkey_data_reg_76));
sg13g2_inv_4 U577 (.A(n1123), .Y(next_addroundkey_round_2));
sg13g2_a21oi_2 U578 (.A1(n1120), .A2(N1537), .B1(n1124), .Y(n1123));
sg13g2_nand3_1 U579 (.A(n1261), .B(n3668), .C(n1260), .Y(next_addroundkey_data_reg_77));
sg13g2_nand3_1 U580 (.A(n1256), .B(n3669), .C(n1255), .Y(next_addroundkey_data_reg_78));
sg13g2_nand3_1 U581 (.A(n1251), .B(n3670), .C(n1250), .Y(next_addroundkey_data_reg_79));
sg13g2_nand3_1 U582 (.A(n1246), .B(n3671), .C(n1245), .Y(next_addroundkey_data_reg_7));
sg13g2_inv_4 U583 (.A(n1127), .Y(n1120));
sg13g2_nand3_1 U584 (.A(n1241), .B(n3672), .C(n1240), .Y(next_addroundkey_data_reg_80));
sg13g2_nand2_2 U585 (.A(addroundkey_round_0), .B(n1129), .Y(n1128));
sg13g2_inv_4 U586 (.A(n1122), .Y(n1129));
sg13g2_nand3_1 U587 (.A(net39311), .B(n1131), .C(n168), .Y(n1122));
sg13g2_nand3_1 U588 (.A(keysched_ready_o), .B(net39311), .C(n168), .Y(n1127));
sg13g2_nand3_1 U589 (.A(n1236), .B(n3673), .C(n1235), .Y(next_addroundkey_data_reg_81));
sg13g2_a21oi_2 U590 (.A1(net24687), .A2(N848), .B1(n1135), .Y(n1133));
sg13g2_nor2_2 U591 (.A(n1136), .B(n4278), .Y(n1135));
sg13g2_a21oi_2 U592 (.A1(net24743), .A2(N1104), .B1(n1139), .Y(n1132));
sg13g2_nor2_2 U593 (.A(n46), .B(n4282), .Y(n1139));
sg13g2_nand3_1 U594 (.A(n1231), .B(n3674), .C(n1230), .Y(next_addroundkey_data_reg_82));
sg13g2_a21oi_2 U595 (.A1(net24687), .A2(N758), .B1(n1142), .Y(n1141));
sg13g2_nor2_2 U596 (.A(n1143), .B(n4278), .Y(n1142));
sg13g2_a21oi_2 U597 (.A1(net24743), .A2(N1014), .B1(n1144), .Y(n1140));
sg13g2_nor2_2 U598 (.A(n136), .B(n4282), .Y(n1144));
sg13g2_nand3_1 U599 (.A(n1226), .B(n3675), .C(n1225), .Y(next_addroundkey_data_reg_83));
sg13g2_a21oi_2 U600 (.A1(net24685), .A2(N759), .B1(n1147), .Y(n1146));
sg13g2_nor2_2 U601 (.A(n1148), .B(n4278), .Y(n1147));
sg13g2_a21oi_2 U602 (.A1(net24743), .A2(N1015), .B1(n1149), .Y(n1145));
sg13g2_nor2_2 U603 (.A(n135), .B(n4282), .Y(n1149));
sg13g2_nand3_1 U604 (.A(n1221), .B(n3677), .C(n1220), .Y(next_addroundkey_data_reg_84));
sg13g2_a21oi_2 U605 (.A1(net24685), .A2(N760), .B1(n1152), .Y(n1151));
sg13g2_nor2_2 U606 (.A(n1153), .B(n4278), .Y(n1152));
sg13g2_a21oi_2 U607 (.A1(net24743), .A2(N1016), .B1(n1154), .Y(n1150));
sg13g2_nor2_2 U608 (.A(n134), .B(n4282), .Y(n1154));
sg13g2_nand3_1 U609 (.A(n1216), .B(n3678), .C(n1215), .Y(next_addroundkey_data_reg_85));
sg13g2_a21oi_2 U610 (.A1(net24687), .A2(N761), .B1(n1157), .Y(n1156));
sg13g2_nor2_2 U611 (.A(n1158), .B(n4278), .Y(n1157));
sg13g2_a21oi_2 U612 (.A1(net24743), .A2(N1017), .B1(n1159), .Y(n1155));
sg13g2_nor2_2 U613 (.A(n133), .B(n4282), .Y(n1159));
sg13g2_nand3_1 U614 (.A(n1211), .B(n3679), .C(n1210), .Y(next_addroundkey_data_reg_86));
sg13g2_a21oi_2 U615 (.A1(net24689), .A2(N762), .B1(n1162), .Y(n1161));
sg13g2_nor2_2 U616 (.A(n1163), .B(n4278), .Y(n1162));
sg13g2_a21oi_2 U617 (.A1(net24743), .A2(N1018), .B1(n1164), .Y(n1160));
sg13g2_nor2_2 U618 (.A(n132), .B(n4282), .Y(n1164));
sg13g2_nand3_1 U619 (.A(n1206), .B(n3680), .C(n1205), .Y(next_addroundkey_data_reg_87));
sg13g2_a21oi_2 U620 (.A1(net24687), .A2(N763), .B1(n1167), .Y(n1166));
sg13g2_nor2_2 U621 (.A(n1168), .B(n4278), .Y(n1167));
sg13g2_a21oi_2 U622 (.A1(net24743), .A2(N1019), .B1(n1169), .Y(n1165));
sg13g2_nor2_2 U623 (.A(n131), .B(n4282), .Y(n1169));
sg13g2_nand3_1 U624 (.A(n1201), .B(n3685), .C(n1200), .Y(next_addroundkey_data_reg_88));
sg13g2_a21oi_2 U625 (.A1(net24689), .A2(N764), .B1(n1172), .Y(n1171));
sg13g2_nor2_2 U626 (.A(n1173), .B(n4278), .Y(n1172));
sg13g2_a21oi_2 U627 (.A1(net24743), .A2(N1020), .B1(n1174), .Y(n1170));
sg13g2_nor2_2 U628 (.A(n130), .B(n4282), .Y(n1174));
sg13g2_nand3_1 U629 (.A(n1196), .B(n3686), .C(n1195), .Y(next_addroundkey_data_reg_89));
sg13g2_a21oi_2 U630 (.A1(net24687), .A2(N765), .B1(n1177), .Y(n1176));
sg13g2_nor2_2 U631 (.A(n1178), .B(n4278), .Y(n1177));
sg13g2_a21oi_2 U632 (.A1(net24743), .A2(N1021), .B1(n1179), .Y(n1175));
sg13g2_nor2_2 U633 (.A(n129), .B(n4282), .Y(n1179));
sg13g2_nand3_1 U634 (.A(n1191), .B(n3687), .C(n1190), .Y(next_addroundkey_data_reg_8));
sg13g2_a21oi_2 U635 (.A1(net24689), .A2(N766), .B1(n1182), .Y(n1181));
sg13g2_nor2_2 U636 (.A(n1183), .B(n4278), .Y(n1182));
sg13g2_a21oi_2 U637 (.A1(net24743), .A2(N1022), .B1(n1184), .Y(n1180));
sg13g2_nor2_2 U638 (.A(n128), .B(n4282), .Y(n1184));
sg13g2_nand3_1 U639 (.A(n1186), .B(n3690), .C(n1185), .Y(next_addroundkey_data_reg_90));
sg13g2_a21oi_2 U640 (.A1(net24689), .A2(N767), .B1(n1187), .Y(n1186));
sg13g2_nor2_2 U641 (.A(n1188), .B(n4278), .Y(n1187));
sg13g2_a21oi_2 U642 (.A1(net24743), .A2(N1023), .B1(n1189), .Y(n1185));
sg13g2_nor2_2 U643 (.A(n127), .B(n4282), .Y(n1189));
sg13g2_nand3_1 U644 (.A(n1181), .B(n3698), .C(n1180), .Y(next_addroundkey_data_reg_91));
sg13g2_a21oi_2 U645 (.A1(net24687), .A2(N849), .B1(n1192), .Y(n1191));
sg13g2_nor2_2 U646 (.A(n1193), .B(n4278), .Y(n1192));
sg13g2_a21oi_2 U647 (.A1(net24743), .A2(N1105), .B1(n1194), .Y(n1190));
sg13g2_nor2_2 U648 (.A(n45), .B(net24601), .Y(n1194));
sg13g2_nand3_1 U649 (.A(n1176), .B(n3709), .C(n1175), .Y(next_addroundkey_data_reg_92));
sg13g2_a21oi_2 U650 (.A1(net24689), .A2(N768), .B1(n1197), .Y(n1196));
sg13g2_nor2_2 U651 (.A(n1198), .B(n4278), .Y(n1197));
sg13g2_a21oi_2 U652 (.A1(net24743), .A2(N1024), .B1(n1199), .Y(n1195));
sg13g2_nor2_2 U653 (.A(n126), .B(net24601), .Y(n1199));
sg13g2_nand3_1 U654 (.A(n1171), .B(n3711), .C(n1170), .Y(next_addroundkey_data_reg_93));
sg13g2_a21oi_2 U655 (.A1(net24685), .A2(N769), .B1(n1202), .Y(n1201));
sg13g2_nor2_2 U656 (.A(n1203), .B(n4278), .Y(n1202));
sg13g2_a21oi_2 U657 (.A1(net24743), .A2(N1025), .B1(n1204), .Y(n1200));
sg13g2_nor2_2 U658 (.A(n125), .B(net24601), .Y(n1204));
sg13g2_nand3_1 U659 (.A(n1166), .B(n3712), .C(n1165), .Y(next_addroundkey_data_reg_94));
sg13g2_a21oi_2 U660 (.A1(net24689), .A2(N770), .B1(n1207), .Y(n1206));
sg13g2_nor2_2 U661 (.A(n1208), .B(n4278), .Y(n1207));
sg13g2_a21oi_2 U662 (.A1(net24743), .A2(N1026), .B1(n1209), .Y(n1205));
sg13g2_nor2_2 U663 (.A(n124), .B(net24601), .Y(n1209));
sg13g2_nand3_1 U664 (.A(n1161), .B(n3713), .C(n1160), .Y(next_addroundkey_data_reg_95));
sg13g2_a21oi_2 U665 (.A1(net24687), .A2(N771), .B1(n1212), .Y(n1211));
sg13g2_nor2_2 U666 (.A(n1213), .B(n4278), .Y(n1212));
sg13g2_a21oi_2 U667 (.A1(net24743), .A2(N1027), .B1(n1214), .Y(n1210));
sg13g2_nor2_2 U668 (.A(n123), .B(net24601), .Y(n1214));
sg13g2_nand3_1 U669 (.A(n1156), .B(n3717), .C(n1155), .Y(next_addroundkey_data_reg_96));
sg13g2_a21oi_2 U670 (.A1(net24689), .A2(N772), .B1(n1217), .Y(n1216));
sg13g2_nor2_2 U671 (.A(n1218), .B(n4278), .Y(n1217));
sg13g2_a21oi_2 U672 (.A1(net24743), .A2(N1028), .B1(n1219), .Y(n1215));
sg13g2_nor2_2 U673 (.A(n122), .B(net24601), .Y(n1219));
sg13g2_nand3_1 U674 (.A(n1151), .B(n3720), .C(n1150), .Y(next_addroundkey_data_reg_97));
sg13g2_a21oi_2 U675 (.A1(net24689), .A2(N773), .B1(n1222), .Y(n1221));
sg13g2_nor2_2 U676 (.A(n1223), .B(n4278), .Y(n1222));
sg13g2_a21oi_2 U677 (.A1(net24743), .A2(N1029), .B1(n1224), .Y(n1220));
sg13g2_nor2_2 U678 (.A(n121), .B(net24601), .Y(n1224));
sg13g2_nand3_1 U679 (.A(n1146), .B(n3723), .C(n1145), .Y(next_addroundkey_data_reg_98));
sg13g2_a21oi_2 U680 (.A1(net24687), .A2(N774), .B1(n1227), .Y(n1226));
sg13g2_nor2_2 U681 (.A(n1228), .B(n4278), .Y(n1227));
sg13g2_a21oi_2 U682 (.A1(net24743), .A2(N1030), .B1(n1229), .Y(n1225));
sg13g2_nor2_2 U683 (.A(n120), .B(net24601), .Y(n1229));
sg13g2_nand3_1 U684 (.A(n1141), .B(n3724), .C(n1140), .Y(next_addroundkey_data_reg_99));
sg13g2_a21oi_2 U685 (.A1(net24685), .A2(N775), .B1(n1232), .Y(n1231));
sg13g2_nor2_2 U686 (.A(n1233), .B(n4278), .Y(n1232));
sg13g2_a21oi_2 U687 (.A1(net24743), .A2(N1031), .B1(n1234), .Y(n1230));
sg13g2_nor2_2 U688 (.A(n119), .B(net24601), .Y(n1234));
sg13g2_nand3_1 U689 (.A(n1133), .B(n3726), .C(n1132), .Y(next_addroundkey_data_reg_9));
sg13g2_a21oi_2 U690 (.A1(net24687), .A2(N776), .B1(n1237), .Y(n1236));
sg13g2_nor2_2 U691 (.A(n1238), .B(n4278), .Y(n1237));
sg13g2_a21oi_2 U692 (.A1(net24743), .A2(N1032), .B1(n1239), .Y(n1235));
sg13g2_nor2_2 U693 (.A(n118), .B(net24601), .Y(n1239));
sg13g2_nand3_1 U694 (.A(n168), .B(n3735), .C(n1128), .Y(next_addroundkey_round_0));
sg13g2_a21oi_2 U695 (.A1(net24685), .A2(N777), .B1(n1242), .Y(n1241));
sg13g2_nor2_2 U696 (.A(n1243), .B(n4278), .Y(n1242));
sg13g2_a21oi_2 U697 (.A1(net24743), .A2(N1033), .B1(n1244), .Y(n1240));
sg13g2_nor2_2 U698 (.A(n117), .B(net24601), .Y(n1244));
sg13g2_nor2_1 U699 (.A(n3693), .B(n3688), .Y(n1));
sg13g2_a21oi_2 U700 (.A1(net24689), .A2(N850), .B1(n1247), .Y(n1246));
sg13g2_nor2_2 U701 (.A(n1248), .B(n4278), .Y(n1247));
sg13g2_a21oi_2 U702 (.A1(net24743), .A2(N1106), .B1(n1249), .Y(n1245));
sg13g2_nor2_2 U703 (.A(n44), .B(net24601), .Y(n1249));
sg13g2_nand2_1 U704 (.A(n1120), .B(n3736), .Y(n3735));
sg13g2_a21oi_2 U705 (.A1(net24685), .A2(N778), .B1(n1252), .Y(n1251));
sg13g2_nor2_2 U706 (.A(n1253), .B(n4278), .Y(n1252));
sg13g2_a21oi_2 U707 (.A1(net24743), .A2(N1034), .B1(n1254), .Y(n1250));
sg13g2_nor2_2 U708 (.A(n116), .B(net24601), .Y(n1254));
sg13g2_or2_1 U709 (.A(n4281), .B(n306), .X(n3726));
sg13g2_a21oi_2 U710 (.A1(net24689), .A2(N779), .B1(n1257), .Y(n1256));
sg13g2_nor2_2 U711 (.A(n1258), .B(n4278), .Y(n1257));
sg13g2_a21oi_2 U712 (.A1(net24743), .A2(N1035), .B1(n1259), .Y(n1255));
sg13g2_nor2_2 U713 (.A(n115), .B(net24601), .Y(n1259));
sg13g2_or2_1 U714 (.A(n4281), .B(n396), .X(n3724));
sg13g2_a21oi_2 U715 (.A1(net24689), .A2(N780), .B1(n1262), .Y(n1261));
sg13g2_nor2_2 U716 (.A(n1263), .B(n4278), .Y(n1262));
sg13g2_a21oi_2 U717 (.A1(net24743), .A2(N1036), .B1(n1264), .Y(n1260));
sg13g2_nor2_2 U718 (.A(n114), .B(net24601), .Y(n1264));
sg13g2_or2_1 U719 (.A(n4281), .B(n395), .X(n3723));
sg13g2_a21oi_2 U720 (.A1(net24685), .A2(N781), .B1(n1267), .Y(n1266));
sg13g2_nor2_2 U721 (.A(n1268), .B(n4278), .Y(n1267));
sg13g2_a21oi_2 U722 (.A1(net24743), .A2(N1037), .B1(n1269), .Y(n1265));
sg13g2_nor2_2 U723 (.A(n113), .B(net24601), .Y(n1269));
sg13g2_or2_1 U724 (.A(n4281), .B(n394), .X(n3720));
sg13g2_a21oi_2 U725 (.A1(net24685), .A2(N782), .B1(n1272), .Y(n1271));
sg13g2_nor2_2 U726 (.A(n1273), .B(n4278), .Y(n1272));
sg13g2_a21oi_2 U727 (.A1(net24743), .A2(N1038), .B1(n1274), .Y(n1270));
sg13g2_nor2_2 U728 (.A(n112), .B(net24601), .Y(n1274));
sg13g2_or2_1 U729 (.A(n4281), .B(n393), .X(n3717));
sg13g2_a21oi_2 U730 (.A1(n1134), .A2(N783), .B1(n1277), .Y(n1276));
sg13g2_nor2_2 U731 (.A(n1278), .B(n4278), .Y(n1277));
sg13g2_a21oi_2 U732 (.A1(net24743), .A2(N1039), .B1(n1279), .Y(n1275));
sg13g2_nor2_2 U733 (.A(n111), .B(net24601), .Y(n1279));
sg13g2_or2_1 U734 (.A(n4281), .B(n392), .X(n3713));
sg13g2_a21oi_2 U735 (.A1(net24687), .A2(N784), .B1(n1282), .Y(n1281));
sg13g2_nor2_2 U736 (.A(n1283), .B(n4278), .Y(n1282));
sg13g2_a21oi_2 U737 (.A1(net24743), .A2(N1040), .B1(n1284), .Y(n1280));
sg13g2_nor2_2 U738 (.A(n110), .B(net24601), .Y(n1284));
sg13g2_or2_1 U739 (.A(n4281), .B(n391), .X(n3712));
sg13g2_a21oi_2 U740 (.A1(n1134), .A2(N785), .B1(n1287), .Y(n1286));
sg13g2_nor2_2 U741 (.A(n1288), .B(n4278), .Y(n1287));
sg13g2_a21oi_2 U742 (.A1(net24743), .A2(N1041), .B1(n1289), .Y(n1285));
sg13g2_nor2_2 U743 (.A(n109), .B(net24601), .Y(n1289));
sg13g2_or2_1 U744 (.A(n4281), .B(n390), .X(n3711));
sg13g2_a21oi_2 U745 (.A1(net24689), .A2(N786), .B1(n1292), .Y(n1291));
sg13g2_nor2_2 U746 (.A(n1293), .B(n4278), .Y(n1292));
sg13g2_a21oi_2 U747 (.A1(net24743), .A2(N1042), .B1(n1294), .Y(n1290));
sg13g2_nor2_2 U748 (.A(n108), .B(n4282), .Y(n1294));
sg13g2_or2_1 U749 (.A(n4281), .B(n389), .X(n3709));
sg13g2_a21oi_2 U750 (.A1(net24689), .A2(N787), .B1(n1297), .Y(n1296));
sg13g2_nor2_2 U751 (.A(n1298), .B(n4278), .Y(n1297));
sg13g2_a21oi_2 U752 (.A1(net24743), .A2(N1043), .B1(n1299), .Y(n1295));
sg13g2_nor2_2 U753 (.A(n107), .B(net24601), .Y(n1299));
sg13g2_or2_1 U754 (.A(n4281), .B(n388), .X(n3698));
sg13g2_a21oi_2 U755 (.A1(n1134), .A2(N851), .B1(n1302), .Y(n1301));
sg13g2_nor2_2 U756 (.A(n1303), .B(n4278), .Y(n1302));
sg13g2_a21oi_2 U757 (.A1(net24743), .A2(N1107), .B1(n1304), .Y(n1300));
sg13g2_nor2_2 U758 (.A(n43), .B(net24601), .Y(n1304));
sg13g2_or2_1 U759 (.A(n4281), .B(n387), .X(n3690));
sg13g2_a21oi_2 U760 (.A1(net24685), .A2(N788), .B1(n1307), .Y(n1306));
sg13g2_nor2_2 U761 (.A(n1308), .B(n4278), .Y(n1307));
sg13g2_a21oi_2 U762 (.A1(net24743), .A2(N1044), .B1(n1309), .Y(n1305));
sg13g2_nor2_2 U763 (.A(n106), .B(net24611), .Y(n1309));
sg13g2_or2_1 U764 (.A(n4281), .B(n305), .X(n3687));
sg13g2_a21oi_2 U765 (.A1(net24689), .A2(N789), .B1(n1312), .Y(n1311));
sg13g2_nor2_2 U766 (.A(n1313), .B(n4278), .Y(n1312));
sg13g2_a21oi_2 U767 (.A1(net24743), .A2(N1045), .B1(n1314), .Y(n1310));
sg13g2_nor2_2 U768 (.A(n105), .B(net24611), .Y(n1314));
sg13g2_or2_1 U769 (.A(n4281), .B(n386), .X(n3686));
sg13g2_a21oi_2 U770 (.A1(net24689), .A2(N790), .B1(n1317), .Y(n1316));
sg13g2_nor2_2 U771 (.A(n1318), .B(n4278), .Y(n1317));
sg13g2_a21oi_2 U772 (.A1(net24743), .A2(N1046), .B1(n1319), .Y(n1315));
sg13g2_nor2_2 U773 (.A(n104), .B(net24611), .Y(n1319));
sg13g2_or2_1 U774 (.A(n4281), .B(n385), .X(n3685));
sg13g2_a21oi_2 U775 (.A1(net24687), .A2(N791), .B1(n1322), .Y(n1321));
sg13g2_nor2_2 U776 (.A(n1323), .B(n4278), .Y(n1322));
sg13g2_a21oi_2 U777 (.A1(net24743), .A2(N1047), .B1(n1324), .Y(n1320));
sg13g2_nor2_2 U778 (.A(n103), .B(net24611), .Y(n1324));
sg13g2_or2_1 U779 (.A(n4281), .B(n384), .X(n3680));
sg13g2_a21oi_2 U780 (.A1(net24685), .A2(N792), .B1(n1327), .Y(n1326));
sg13g2_nor2_2 U781 (.A(n1328), .B(n4278), .Y(n1327));
sg13g2_a21oi_2 U782 (.A1(net24743), .A2(N1048), .B1(n1329), .Y(n1325));
sg13g2_nor2_2 U783 (.A(n102), .B(n4282), .Y(n1329));
sg13g2_or2_1 U784 (.A(n4281), .B(n383), .X(n3679));
sg13g2_a21oi_2 U785 (.A1(net24685), .A2(N793), .B1(n1332), .Y(n1331));
sg13g2_nor2_2 U786 (.A(n1333), .B(n4278), .Y(n1332));
sg13g2_a21oi_2 U787 (.A1(net24743), .A2(N1049), .B1(n1334), .Y(n1330));
sg13g2_nor2_2 U788 (.A(n101), .B(n4282), .Y(n1334));
sg13g2_or2_1 U789 (.A(n4281), .B(n382), .X(n3678));
sg13g2_a21oi_2 U790 (.A1(net24687), .A2(N794), .B1(n1337), .Y(n1336));
sg13g2_nor2_2 U791 (.A(n1338), .B(n4278), .Y(n1337));
sg13g2_a21oi_2 U792 (.A1(net24743), .A2(N1050), .B1(n1339), .Y(n1335));
sg13g2_nor2_2 U793 (.A(n100), .B(n4282), .Y(n1339));
sg13g2_or2_1 U794 (.A(n4281), .B(n381), .X(n3677));
sg13g2_a21oi_2 U795 (.A1(net24685), .A2(N795), .B1(n1342), .Y(n1341));
sg13g2_nor2_2 U796 (.A(n1343), .B(n4278), .Y(n1342));
sg13g2_a21oi_2 U797 (.A1(net24743), .A2(N1051), .B1(n1344), .Y(n1340));
sg13g2_nor2_2 U798 (.A(n99), .B(net24611), .Y(n1344));
sg13g2_or2_1 U799 (.A(n4281), .B(n380), .X(n3675));
sg13g2_a21oi_2 U800 (.A1(net24689), .A2(N796), .B1(n1347), .Y(n1346));
sg13g2_nor2_2 U801 (.A(n1348), .B(n4278), .Y(n1347));
sg13g2_a21oi_2 U802 (.A1(net24743), .A2(N1052), .B1(n1349), .Y(n1345));
sg13g2_nor2_2 U803 (.A(n98), .B(n4282), .Y(n1349));
sg13g2_or2_1 U804 (.A(n4281), .B(n379), .X(n3674));
sg13g2_a21oi_2 U805 (.A1(net24687), .A2(N797), .B1(n1352), .Y(n1351));
sg13g2_nor2_2 U806 (.A(n1353), .B(n4278), .Y(n1352));
sg13g2_a21oi_2 U807 (.A1(net24743), .A2(N1053), .B1(n1354), .Y(n1350));
sg13g2_nor2_2 U808 (.A(n97), .B(net24611), .Y(n1354));
sg13g2_or2_1 U809 (.A(n4281), .B(n378), .X(n3673));
sg13g2_a21oi_2 U810 (.A1(net24685), .A2(N852), .B1(n1357), .Y(n1356));
sg13g2_nor2_2 U811 (.A(n1358), .B(n4278), .Y(n1357));
sg13g2_a21oi_2 U812 (.A1(net24743), .A2(N1108), .B1(n1359), .Y(n1355));
sg13g2_nor2_2 U813 (.A(n42), .B(net24611), .Y(n1359));
sg13g2_or2_1 U814 (.A(n4281), .B(n377), .X(n3672));
sg13g2_a21oi_2 U815 (.A1(net24685), .A2(N798), .B1(n1362), .Y(n1361));
sg13g2_nor2_2 U816 (.A(n1363), .B(n4278), .Y(n1362));
sg13g2_a21oi_2 U817 (.A1(net24743), .A2(N1054), .B1(n1364), .Y(n1360));
sg13g2_nor2_2 U818 (.A(n96), .B(net24611), .Y(n1364));
sg13g2_or2_1 U819 (.A(n4281), .B(n304), .X(n3671));
sg13g2_a21oi_2 U820 (.A1(net24689), .A2(N799), .B1(n1367), .Y(n1366));
sg13g2_nor2_2 U821 (.A(n1368), .B(n4278), .Y(n1367));
sg13g2_a21oi_2 U822 (.A1(net24743), .A2(N1055), .B1(n1369), .Y(n1365));
sg13g2_nor2_2 U823 (.A(n95), .B(n4282), .Y(n1369));
sg13g2_or2_1 U824 (.A(n4281), .B(n376), .X(n3670));
sg13g2_a21oi_2 U825 (.A1(net24689), .A2(N800), .B1(n1372), .Y(n1371));
sg13g2_nor2_2 U826 (.A(n1373), .B(n4278), .Y(n1372));
sg13g2_a21oi_2 U827 (.A1(net24743), .A2(N1056), .B1(n1374), .Y(n1370));
sg13g2_nor2_2 U828 (.A(n94), .B(n4282), .Y(n1374));
sg13g2_or2_1 U829 (.A(n4281), .B(n375), .X(n3669));
sg13g2_a21oi_2 U830 (.A1(net24685), .A2(N801), .B1(n1377), .Y(n1376));
sg13g2_nor2_2 U831 (.A(n1378), .B(n4278), .Y(n1377));
sg13g2_a21oi_2 U832 (.A1(net24743), .A2(N1057), .B1(n1379), .Y(n1375));
sg13g2_nor2_2 U833 (.A(n93), .B(n4282), .Y(n1379));
sg13g2_or2_1 U834 (.A(n4281), .B(n374), .X(n3668));
sg13g2_a21oi_2 U835 (.A1(net24687), .A2(N802), .B1(n1382), .Y(n1381));
sg13g2_nor2_2 U836 (.A(n1383), .B(n4278), .Y(n1382));
sg13g2_a21oi_2 U837 (.A1(net24743), .A2(N1058), .B1(n1384), .Y(n1380));
sg13g2_nor2_2 U838 (.A(n92), .B(net24611), .Y(n1384));
sg13g2_or2_1 U839 (.A(n4281), .B(n373), .X(n3667));
sg13g2_a21oi_2 U840 (.A1(net24685), .A2(N803), .B1(n1387), .Y(n1386));
sg13g2_nor2_2 U841 (.A(n1388), .B(n4278), .Y(n1387));
sg13g2_a21oi_2 U842 (.A1(net24743), .A2(N1059), .B1(n1389), .Y(n1385));
sg13g2_nor2_2 U843 (.A(n91), .B(n4282), .Y(n1389));
sg13g2_or2_1 U844 (.A(n4281), .B(n372), .X(n3666));
sg13g2_a21oi_2 U845 (.A1(n1134), .A2(N804), .B1(n1392), .Y(n1391));
sg13g2_nor2_2 U846 (.A(n1393), .B(n4278), .Y(n1392));
sg13g2_a21oi_2 U847 (.A1(net24743), .A2(N1060), .B1(n1394), .Y(n1390));
sg13g2_nor2_2 U848 (.A(n90), .B(n4282), .Y(n1394));
sg13g2_or2_1 U849 (.A(n4281), .B(n371), .X(n3665));
sg13g2_a21oi_2 U850 (.A1(net24685), .A2(N805), .B1(n1397), .Y(n1396));
sg13g2_nor2_2 U851 (.A(n1398), .B(n4278), .Y(n1397));
sg13g2_a21oi_2 U852 (.A1(net24743), .A2(N1061), .B1(n1399), .Y(n1395));
sg13g2_nor2_2 U853 (.A(n89), .B(n4282), .Y(n1399));
sg13g2_or2_1 U854 (.A(n4281), .B(n370), .X(n3664));
sg13g2_a21oi_2 U855 (.A1(n1134), .A2(N806), .B1(n1402), .Y(n1401));
sg13g2_nor2_2 U856 (.A(n1403), .B(n4278), .Y(n1402));
sg13g2_a21oi_2 U857 (.A1(net24743), .A2(N1062), .B1(n1404), .Y(n1400));
sg13g2_nor2_2 U858 (.A(n88), .B(n4282), .Y(n1404));
sg13g2_or2_1 U859 (.A(n4281), .B(n369), .X(n3663));
sg13g2_a21oi_2 U860 (.A1(net24687), .A2(N807), .B1(n1407), .Y(n1406));
sg13g2_nor2_2 U861 (.A(n1408), .B(n4278), .Y(n1407));
sg13g2_a21oi_2 U862 (.A1(net24743), .A2(N1063), .B1(n1409), .Y(n1405));
sg13g2_nor2_2 U863 (.A(n87), .B(n4282), .Y(n1409));
sg13g2_or2_1 U864 (.A(n4281), .B(n368), .X(n3662));
sg13g2_a21oi_2 U865 (.A1(net24687), .A2(N853), .B1(n1412), .Y(n1411));
sg13g2_nor2_2 U866 (.A(n1413), .B(n4278), .Y(n1412));
sg13g2_a21oi_2 U867 (.A1(net24743), .A2(N1109), .B1(n1414), .Y(n1410));
sg13g2_nor2_2 U868 (.A(n41), .B(n4282), .Y(n1414));
sg13g2_or2_1 U869 (.A(n4281), .B(n367), .X(n3661));
sg13g2_a21oi_2 U870 (.A1(net24689), .A2(N808), .B1(n1417), .Y(n1416));
sg13g2_nor2_2 U871 (.A(n1418), .B(n4278), .Y(n1417));
sg13g2_a21oi_2 U872 (.A1(net24743), .A2(N1064), .B1(n1419), .Y(n1415));
sg13g2_nor2_2 U873 (.A(n86), .B(net24611), .Y(n1419));
sg13g2_or2_1 U874 (.A(n4281), .B(n303), .X(n3660));
sg13g2_a21oi_2 U875 (.A1(net24689), .A2(N809), .B1(n1422), .Y(n1421));
sg13g2_nor2_2 U876 (.A(n1423), .B(n4278), .Y(n1422));
sg13g2_a21oi_2 U877 (.A1(net24743), .A2(N1065), .B1(n1424), .Y(n1420));
sg13g2_nor2_2 U878 (.A(n85), .B(net24611), .Y(n1424));
sg13g2_or2_1 U879 (.A(n4281), .B(n366), .X(n3659));
sg13g2_a21oi_2 U880 (.A1(net24687), .A2(N810), .B1(n1427), .Y(n1426));
sg13g2_nor2_2 U881 (.A(n1428), .B(n4278), .Y(n1427));
sg13g2_a21oi_2 U882 (.A1(net24743), .A2(N1066), .B1(n1429), .Y(n1425));
sg13g2_nor2_2 U883 (.A(n84), .B(n4282), .Y(n1429));
sg13g2_or2_1 U884 (.A(n4281), .B(n365), .X(n3658));
sg13g2_a21oi_2 U885 (.A1(net24687), .A2(N811), .B1(n1432), .Y(n1431));
sg13g2_nor2_2 U886 (.A(n1433), .B(n4278), .Y(n1432));
sg13g2_a21oi_2 U887 (.A1(net24743), .A2(N1067), .B1(n1434), .Y(n1430));
sg13g2_nor2_2 U888 (.A(n83), .B(net24601), .Y(n1434));
sg13g2_or2_1 U889 (.A(n4281), .B(n364), .X(n3524));
sg13g2_a21oi_2 U890 (.A1(net24689), .A2(N812), .B1(n1437), .Y(n1436));
sg13g2_nor2_2 U891 (.A(n1438), .B(n4278), .Y(n1437));
sg13g2_a21oi_2 U892 (.A1(net24743), .A2(N1068), .B1(n1439), .Y(n1435));
sg13g2_nor2_2 U893 (.A(n82), .B(n4282), .Y(n1439));
sg13g2_or2_1 U894 (.A(n4281), .B(n363), .X(n2240));
sg13g2_a21oi_2 U895 (.A1(net24685), .A2(N813), .B1(n1442), .Y(n1441));
sg13g2_nor2_2 U896 (.A(n1443), .B(n4278), .Y(n1442));
sg13g2_a21oi_2 U897 (.A1(net24743), .A2(N1069), .B1(n1444), .Y(n1440));
sg13g2_nor2_2 U898 (.A(n81), .B(net24611), .Y(n1444));
sg13g2_or2_1 U899 (.A(n4281), .B(n362), .X(n2239));
sg13g2_a21oi_2 U900 (.A1(net24687), .A2(N814), .B1(n1447), .Y(n1446));
sg13g2_nor2_2 U901 (.A(n1448), .B(n4278), .Y(n1447));
sg13g2_a21oi_2 U902 (.A1(net24743), .A2(N1070), .B1(n1449), .Y(n1445));
sg13g2_nor2_2 U903 (.A(n80), .B(n4282), .Y(n1449));
sg13g2_or2_1 U904 (.A(n4281), .B(n361), .X(n2238));
sg13g2_a21oi_2 U905 (.A1(net24689), .A2(N815), .B1(n1452), .Y(n1451));
sg13g2_nor2_2 U906 (.A(n1453), .B(n4278), .Y(n1452));
sg13g2_a21oi_2 U907 (.A1(net24743), .A2(N1071), .B1(n1454), .Y(n1450));
sg13g2_nor2_2 U908 (.A(n79), .B(n4282), .Y(n1454));
sg13g2_or2_1 U909 (.A(n4281), .B(n360), .X(n2237));
sg13g2_a21oi_2 U910 (.A1(n1134), .A2(N816), .B1(n1457), .Y(n1456));
sg13g2_nor2_2 U911 (.A(n1458), .B(n4278), .Y(n1457));
sg13g2_a21oi_2 U912 (.A1(net24743), .A2(N1072), .B1(n1459), .Y(n1455));
sg13g2_nor2_2 U913 (.A(n78), .B(net24601), .Y(n1459));
sg13g2_or2_1 U914 (.A(n4281), .B(n359), .X(n2236));
sg13g2_a21oi_2 U915 (.A1(net24689), .A2(N817), .B1(n1462), .Y(n1461));
sg13g2_nor2_2 U916 (.A(n1463), .B(n4278), .Y(n1462));
sg13g2_a21oi_2 U917 (.A1(net24743), .A2(N1073), .B1(n1464), .Y(n1460));
sg13g2_nor2_2 U918 (.A(n77), .B(n4282), .Y(n1464));
sg13g2_or2_1 U919 (.A(n4281), .B(n358), .X(n2173));
sg13g2_a21oi_2 U920 (.A1(net24685), .A2(N854), .B1(n1467), .Y(n1466));
sg13g2_nor2_2 U921 (.A(n1468), .B(n4278), .Y(n1467));
sg13g2_a21oi_2 U922 (.A1(net24743), .A2(N1110), .B1(n1469), .Y(n1465));
sg13g2_nor2_2 U923 (.A(n40), .B(n4282), .Y(n1469));
sg13g2_or2_1 U924 (.A(n4281), .B(n357), .X(n1916));
sg13g2_or2_1 U925 (.A(n4281), .B(n302), .X(n1915));
sg13g2_nor2_2 U926 (.A(n1473), .B(n4278), .Y(n1472));
sg13g2_a21oi_2 U927 (.A1(net24743), .A2(N1074), .B1(n1474), .Y(n1470));
sg13g2_nor2_2 U928 (.A(n76), .B(n4282), .Y(n1474));
sg13g2_or2_1 U929 (.A(n4281), .B(n356), .X(n1908));
sg13g2_a21oi_2 U930 (.A1(net24689), .A2(N819), .B1(n1477), .Y(n1476));
sg13g2_nor2_2 U931 (.A(n1478), .B(n4278), .Y(n1477));
sg13g2_a21oi_2 U932 (.A1(net24743), .A2(N1075), .B1(n1479), .Y(n1475));
sg13g2_nor2_2 U933 (.A(n75), .B(n4282), .Y(n1479));
sg13g2_or2_1 U934 (.A(n4281), .B(n355), .X(n1906));
sg13g2_a21oi_2 U935 (.A1(net24687), .A2(N820), .B1(n1482), .Y(n1481));
sg13g2_nor2_2 U936 (.A(n1483), .B(n4278), .Y(n1482));
sg13g2_a21oi_2 U937 (.A1(net24743), .A2(N1076), .B1(n1484), .Y(n1480));
sg13g2_nor2_2 U938 (.A(n74), .B(n4282), .Y(n1484));
sg13g2_or2_1 U939 (.A(n4281), .B(n354), .X(n1138));
sg13g2_a21oi_2 U940 (.A1(net24687), .A2(N821), .B1(n1487), .Y(n1486));
sg13g2_nor2_2 U941 (.A(n1488), .B(n4278), .Y(n1487));
sg13g2_a21oi_2 U942 (.A1(net24743), .A2(N1077), .B1(n1489), .Y(n1485));
sg13g2_nor2_2 U943 (.A(n73), .B(n4282), .Y(n1489));
sg13g2_or2_1 U944 (.A(n4281), .B(n353), .X(n1137));
sg13g2_a21oi_2 U945 (.A1(net24689), .A2(N822), .B1(n1492), .Y(n1491));
sg13g2_nor2_2 U946 (.A(n1493), .B(n4278), .Y(n1492));
sg13g2_a21oi_2 U947 (.A1(net24743), .A2(N1078), .B1(n1494), .Y(n1490));
sg13g2_nor2_2 U948 (.A(n72), .B(n4282), .Y(n1494));
sg13g2_or2_1 U949 (.A(n4281), .B(n352), .X(n1130));
sg13g2_a21oi_2 U950 (.A1(net24687), .A2(N823), .B1(n1497), .Y(n1496));
sg13g2_nor2_2 U951 (.A(n1498), .B(n4278), .Y(n1497));
sg13g2_a21oi_2 U952 (.A1(net24743), .A2(N1079), .B1(n1499), .Y(n1495));
sg13g2_nor2_2 U953 (.A(n71), .B(n4282), .Y(n1499));
sg13g2_or2_1 U954 (.A(n4281), .B(n351), .X(n1125));
sg13g2_a21oi_2 U955 (.A1(net24689), .A2(N824), .B1(n1502), .Y(n1501));
sg13g2_nor2_2 U956 (.A(n1503), .B(n4278), .Y(n1502));
sg13g2_a21oi_2 U957 (.A1(net24743), .A2(N1080), .B1(n1504), .Y(n1500));
sg13g2_nor2_2 U958 (.A(n70), .B(n4282), .Y(n1504));
sg13g2_or2_1 U959 (.A(n4281), .B(n350), .X(n1114));
sg13g2_a21oi_2 U960 (.A1(net24685), .A2(N825), .B1(n1507), .Y(n1506));
sg13g2_nor2_2 U961 (.A(n1508), .B(n4278), .Y(n1507));
sg13g2_a21oi_2 U962 (.A1(net24743), .A2(N1081), .B1(n1509), .Y(n1505));
sg13g2_nor2_2 U963 (.A(n69), .B(n4282), .Y(n1509));
sg13g2_or2_1 U964 (.A(n4281), .B(n349), .X(n1113));
sg13g2_a21oi_2 U965 (.A1(net24685), .A2(N826), .B1(n1512), .Y(n1511));
sg13g2_nor2_2 U966 (.A(n1513), .B(n4278), .Y(n1512));
sg13g2_a21oi_2 U967 (.A1(net24743), .A2(N1082), .B1(n1514), .Y(n1510));
sg13g2_nor2_2 U968 (.A(n68), .B(n4282), .Y(n1514));
sg13g2_or2_1 U969 (.A(n4281), .B(n348), .X(n1112));
sg13g2_a21oi_2 U970 (.A1(net24685), .A2(N827), .B1(n1517), .Y(n1516));
sg13g2_nor2_2 U971 (.A(n1518), .B(n4278), .Y(n1517));
sg13g2_a21oi_2 U972 (.A1(net24743), .A2(N1083), .B1(n1519), .Y(n1515));
sg13g2_nor2_2 U973 (.A(n67), .B(n4282), .Y(n1519));
sg13g2_or2_1 U974 (.A(n4281), .B(n347), .X(n1111));
sg13g2_a21oi_2 U975 (.A1(net24687), .A2(N855), .B1(n1522), .Y(n1521));
sg13g2_nor2_2 U976 (.A(n1523), .B(n4278), .Y(n1522));
sg13g2_a21oi_2 U977 (.A1(net24743), .A2(N1111), .B1(n1524), .Y(n1520));
sg13g2_nor2_2 U978 (.A(n39), .B(net24611), .Y(n1524));
sg13g2_or2_1 U979 (.A(n4281), .B(n301), .X(n1110));
sg13g2_a21oi_2 U980 (.A1(net24685), .A2(N828), .B1(n1527), .Y(n1526));
sg13g2_nor2_2 U981 (.A(n1528), .B(n4278), .Y(n1527));
sg13g2_a21oi_2 U982 (.A1(net24743), .A2(N1084), .B1(n1529), .Y(n1525));
sg13g2_nor2_2 U983 (.A(n66), .B(net24611), .Y(n1529));
sg13g2_or2_1 U984 (.A(n4281), .B(n346), .X(n854));
sg13g2_a21oi_2 U985 (.A1(net24685), .A2(N829), .B1(n1532), .Y(n1531));
sg13g2_nor2_2 U986 (.A(n1533), .B(n4278), .Y(n1532));
sg13g2_a21oi_2 U987 (.A1(net24743), .A2(N1085), .B1(n1534), .Y(n1530));
sg13g2_nor2_2 U988 (.A(n65), .B(net24611), .Y(n1534));
sg13g2_or2_1 U989 (.A(n4281), .B(n345), .X(n842));
sg13g2_a21oi_2 U990 (.A1(net24689), .A2(N830), .B1(n1537), .Y(n1536));
sg13g2_nor2_2 U991 (.A(n1538), .B(n4278), .Y(n1537));
sg13g2_a21oi_2 U992 (.A1(net24743), .A2(N1086), .B1(n1539), .Y(n1535));
sg13g2_nor2_2 U993 (.A(n64), .B(net24611), .Y(n1539));
sg13g2_or2_1 U994 (.A(n4281), .B(n344), .X(n833));
sg13g2_a21oi_2 U995 (.A1(net24689), .A2(N831), .B1(n1542), .Y(n1541));
sg13g2_nor2_2 U996 (.A(n1543), .B(n4278), .Y(n1542));
sg13g2_a21oi_2 U997 (.A1(net24743), .A2(N1087), .B1(n1544), .Y(n1540));
sg13g2_nor2_2 U998 (.A(n63), .B(net24611), .Y(n1544));
sg13g2_or2_1 U999 (.A(n4281), .B(n343), .X(n831));
sg13g2_a21oi_2 U1000 (.A1(net24687), .A2(N832), .B1(n1547), .Y(n1546));
sg13g2_nor2_2 U1001 (.A(n1548), .B(n4278), .Y(n1547));
sg13g2_a21oi_2 U1002 (.A1(net24743), .A2(N1088), .B1(n1549), .Y(n1545));
sg13g2_nor2_2 U1003 (.A(n62), .B(net24611), .Y(n1549));
sg13g2_or2_1 U1004 (.A(n4281), .B(n342), .X(n829));
sg13g2_a21oi_2 U1005 (.A1(n1134), .A2(N833), .B1(n1552), .Y(n1551));
sg13g2_nor2_2 U1006 (.A(n1553), .B(n4278), .Y(n1552));
sg13g2_a21oi_2 U1007 (.A1(net24743), .A2(N1089), .B1(n1554), .Y(n1550));
sg13g2_nor2_2 U1008 (.A(n61), .B(net24611), .Y(n1554));
sg13g2_or2_1 U1009 (.A(n4281), .B(n341), .X(n827));
sg13g2_a21oi_2 U1010 (.A1(net24685), .A2(N834), .B1(n1557), .Y(n1556));
sg13g2_nor2_2 U1011 (.A(n1558), .B(n4278), .Y(n1557));
sg13g2_a21oi_2 U1012 (.A1(net24743), .A2(N1090), .B1(n1559), .Y(n1555));
sg13g2_nor2_2 U1013 (.A(n60), .B(net24611), .Y(n1559));
sg13g2_or2_1 U1014 (.A(n4281), .B(n340), .X(n825));
sg13g2_a21oi_2 U1015 (.A1(n1134), .A2(N835), .B1(n1562), .Y(n1561));
sg13g2_nor2_2 U1016 (.A(n1563), .B(n4278), .Y(n1562));
sg13g2_a21oi_2 U1017 (.A1(net24743), .A2(N1091), .B1(n1564), .Y(n1560));
sg13g2_nor2_2 U1018 (.A(n59), .B(net24611), .Y(n1564));
sg13g2_or2_1 U1019 (.A(n4281), .B(n339), .X(n823));
sg13g2_a21oi_2 U1020 (.A1(net24685), .A2(N836), .B1(n1567), .Y(n1566));
sg13g2_nor2_2 U1021 (.A(n1568), .B(n4278), .Y(n1567));
sg13g2_a21oi_2 U1022 (.A1(net24743), .A2(N1092), .B1(n1569), .Y(n1565));
sg13g2_nor2_2 U1023 (.A(n58), .B(net24611), .Y(n1569));
sg13g2_or2_1 U1024 (.A(n4281), .B(n338), .X(n821));
sg13g2_a21oi_2 U1025 (.A1(net24689), .A2(N837), .B1(n1572), .Y(n1571));
sg13g2_nor2_2 U1026 (.A(n1573), .B(n4278), .Y(n1572));
sg13g2_a21oi_2 U1027 (.A1(net24743), .A2(N1093), .B1(n1574), .Y(n1570));
sg13g2_nor2_2 U1028 (.A(n57), .B(net24611), .Y(n1574));
sg13g2_or2_1 U1029 (.A(n4281), .B(n337), .X(n819));
sg13g2_a21oi_2 U1030 (.A1(net24687), .A2(N856), .B1(n1577), .Y(n1576));
sg13g2_nor2_2 U1031 (.A(n1578), .B(n4278), .Y(n1577));
sg13g2_a21oi_2 U1032 (.A1(net24743), .A2(N1112), .B1(n1579), .Y(n1575));
sg13g2_nor2_2 U1033 (.A(n38), .B(n4282), .Y(n1579));
sg13g2_or2_1 U1034 (.A(n4281), .B(n300), .X(n817));
sg13g2_a21oi_2 U1035 (.A1(n1134), .A2(N838), .B1(n1582), .Y(n1581));
sg13g2_nor2_2 U1036 (.A(n1583), .B(n4278), .Y(n1582));
sg13g2_a21oi_2 U1037 (.A1(net24743), .A2(N1094), .B1(n1584), .Y(n1580));
sg13g2_nor2_2 U1038 (.A(n56), .B(n4282), .Y(n1584));
sg13g2_or2_1 U1039 (.A(n4281), .B(n336), .X(n816));
sg13g2_a21oi_2 U1040 (.A1(net24689), .A2(N839), .B1(n1587), .Y(n1586));
sg13g2_nor2_2 U1041 (.A(n1588), .B(n4278), .Y(n1587));
sg13g2_a21oi_2 U1042 (.A1(net24743), .A2(N1095), .B1(n1589), .Y(n1585));
sg13g2_nor2_2 U1043 (.A(n55), .B(n4282), .Y(n1589));
sg13g2_or2_1 U1044 (.A(n4281), .B(n335), .X(n556));
sg13g2_a21oi_2 U1045 (.A1(n1134), .A2(N840), .B1(n1592), .Y(n1591));
sg13g2_nor2_2 U1046 (.A(n1593), .B(n4278), .Y(n1592));
sg13g2_a21oi_2 U1047 (.A1(net24743), .A2(N1096), .B1(n1594), .Y(n1590));
sg13g2_nor2_2 U1048 (.A(n54), .B(net24611), .Y(n1594));
sg13g2_or2_1 U1049 (.A(n4281), .B(n334), .X(n548));
sg13g2_a21oi_2 U1050 (.A1(net24685), .A2(N841), .B1(n1597), .Y(n1596));
sg13g2_nor2_2 U1051 (.A(n1598), .B(n4278), .Y(n1597));
sg13g2_a21oi_2 U1052 (.A1(net24743), .A2(N1097), .B1(n1599), .Y(n1595));
sg13g2_nor2_2 U1053 (.A(n53), .B(n4282), .Y(n1599));
sg13g2_or2_1 U1054 (.A(n4281), .B(n333), .X(n547));
sg13g2_a21oi_2 U1055 (.A1(net24689), .A2(N842), .B1(n1602), .Y(n1601));
sg13g2_nor2_2 U1056 (.A(n1603), .B(n4278), .Y(n1602));
sg13g2_a21oi_2 U1057 (.A1(net24743), .A2(N1098), .B1(n1604), .Y(n1600));
sg13g2_nor2_2 U1058 (.A(n52), .B(n4282), .Y(n1604));
sg13g2_or2_1 U1059 (.A(n4281), .B(n332), .X(n546));
sg13g2_a21oi_2 U1060 (.A1(net24687), .A2(N843), .B1(n1607), .Y(n1606));
sg13g2_nor2_2 U1061 (.A(n1608), .B(n4278), .Y(n1607));
sg13g2_a21oi_2 U1062 (.A1(net24743), .A2(N1099), .B1(n1609), .Y(n1605));
sg13g2_nor2_2 U1063 (.A(n51), .B(n4282), .Y(n1609));
sg13g2_or2_1 U1064 (.A(n4281), .B(n331), .X(n545));
sg13g2_a21oi_2 U1065 (.A1(net24685), .A2(N844), .B1(n1612), .Y(n1611));
sg13g2_nor2_2 U1066 (.A(n1613), .B(n4278), .Y(n1612));
sg13g2_a21oi_2 U1067 (.A1(net24743), .A2(N1100), .B1(n1614), .Y(n1610));
sg13g2_nor2_2 U1068 (.A(n50), .B(n4282), .Y(n1614));
sg13g2_or2_1 U1069 (.A(n4281), .B(n330), .X(n544));
sg13g2_a21oi_2 U1070 (.A1(net24689), .A2(N845), .B1(n1617), .Y(n1616));
sg13g2_nor2_2 U1071 (.A(n1618), .B(n4278), .Y(n1617));
sg13g2_a21oi_2 U1072 (.A1(net24743), .A2(N1101), .B1(n1619), .Y(n1615));
sg13g2_nor2_2 U1073 (.A(n49), .B(n4282), .Y(n1619));
sg13g2_or2_1 U1074 (.A(n4281), .B(n329), .X(n543));
sg13g2_a21oi_2 U1075 (.A1(net24687), .A2(N730), .B1(n1622), .Y(n1621));
sg13g2_nor2_2 U1076 (.A(n1623), .B(n4278), .Y(n1622));
sg13g2_a21oi_2 U1077 (.A1(net24743), .A2(N986), .B1(n1624), .Y(n1620));
sg13g2_nor2_2 U1078 (.A(n164), .B(n4282), .Y(n1624));
sg13g2_or2_1 U1079 (.A(n4281), .B(n328), .X(n542));
sg13g2_a21oi_2 U1080 (.A1(net24687), .A2(N731), .B1(n1627), .Y(n1626));
sg13g2_nor2_2 U1081 (.A(n1628), .B(n4278), .Y(n1627));
sg13g2_a21oi_2 U1082 (.A1(net24743), .A2(N987), .B1(n1629), .Y(n1625));
sg13g2_nor2_2 U1083 (.A(n163), .B(n4282), .Y(n1629));
sg13g2_or2_1 U1084 (.A(n4281), .B(n327), .X(n541));
sg13g2_a21oi_2 U1085 (.A1(net24689), .A2(N732), .B1(n1632), .Y(n1631));
sg13g2_nor2_2 U1086 (.A(n1633), .B(n4278), .Y(n1632));
sg13g2_a21oi_2 U1087 (.A1(net24743), .A2(N988), .B1(n1634), .Y(n1630));
sg13g2_nor2_2 U1088 (.A(n162), .B(n4282), .Y(n1634));
sg13g2_or2_1 U1089 (.A(n4281), .B(n299), .X(n540));
sg13g2_a21oi_2 U1090 (.A1(net24685), .A2(N733), .B1(n1637), .Y(n1636));
sg13g2_nor2_2 U1091 (.A(n1638), .B(n4278), .Y(n1637));
sg13g2_a21oi_2 U1092 (.A1(net24743), .A2(N989), .B1(n1639), .Y(n1635));
sg13g2_nor2_2 U1093 (.A(n161), .B(n4282), .Y(n1639));
sg13g2_or2_1 U1094 (.A(n4281), .B(n326), .X(n539));
sg13g2_a21oi_2 U1095 (.A1(net24687), .A2(N734), .B1(n1642), .Y(n1641));
sg13g2_nor2_2 U1096 (.A(n1643), .B(n4278), .Y(n1642));
sg13g2_a21oi_2 U1097 (.A1(net24743), .A2(N990), .B1(n1644), .Y(n1640));
sg13g2_nor2_2 U1098 (.A(n160), .B(n4282), .Y(n1644));
sg13g2_or2_1 U1099 (.A(n4281), .B(n325), .X(n538));
sg13g2_a21oi_2 U1100 (.A1(net24685), .A2(N735), .B1(n1647), .Y(n1646));
sg13g2_nor2_2 U1101 (.A(n1648), .B(n4278), .Y(n1647));
sg13g2_a21oi_2 U1102 (.A1(net24743), .A2(N991), .B1(n1649), .Y(n1645));
sg13g2_nor2_2 U1103 (.A(n159), .B(n4282), .Y(n1649));
sg13g2_or2_1 U1104 (.A(n4281), .B(n324), .X(n537));
sg13g2_a21oi_2 U1105 (.A1(net24687), .A2(N736), .B1(n1652), .Y(n1651));
sg13g2_nor2_2 U1106 (.A(n1653), .B(n4278), .Y(n1652));
sg13g2_a21oi_2 U1107 (.A1(net24743), .A2(N992), .B1(n1654), .Y(n1650));
sg13g2_nor2_2 U1108 (.A(n158), .B(n4282), .Y(n1654));
sg13g2_or2_1 U1109 (.A(n4281), .B(n323), .X(n536));
sg13g2_a21oi_2 U1110 (.A1(net24689), .A2(N737), .B1(n1657), .Y(n1656));
sg13g2_nor2_2 U1111 (.A(n1658), .B(n4278), .Y(n1657));
sg13g2_a21oi_2 U1112 (.A1(net24743), .A2(N993), .B1(n1659), .Y(n1655));
sg13g2_nor2_2 U1113 (.A(n157), .B(n4282), .Y(n1659));
sg13g2_or2_1 U1114 (.A(n4281), .B(n322), .X(n535));
sg13g2_a21oi_2 U1115 (.A1(n1134), .A2(N846), .B1(n1662), .Y(n1661));
sg13g2_nor2_2 U1116 (.A(n1663), .B(n4278), .Y(n1662));
sg13g2_a21oi_2 U1117 (.A1(net24743), .A2(N1102), .B1(n1664), .Y(n1660));
sg13g2_nor2_2 U1118 (.A(n48), .B(n4282), .Y(n1664));
sg13g2_or2_1 U1119 (.A(n4281), .B(n321), .X(n534));
sg13g2_a21oi_2 U1120 (.A1(net24687), .A2(N738), .B1(n1667), .Y(n1666));
sg13g2_nor2_2 U1121 (.A(n1668), .B(n4278), .Y(n1667));
sg13g2_a21oi_2 U1122 (.A1(net24743), .A2(N994), .B1(n1669), .Y(n1665));
sg13g2_nor2_2 U1123 (.A(n156), .B(n4282), .Y(n1669));
sg13g2_or2_1 U1124 (.A(n4281), .B(n320), .X(n533));
sg13g2_a21oi_2 U1125 (.A1(net24689), .A2(N739), .B1(n1672), .Y(n1671));
sg13g2_nor2_2 U1126 (.A(n1673), .B(n4278), .Y(n1672));
sg13g2_a21oi_2 U1127 (.A1(net24743), .A2(N995), .B1(n1674), .Y(n1670));
sg13g2_nor2_2 U1128 (.A(n155), .B(n4282), .Y(n1674));
sg13g2_or2_1 U1129 (.A(n4281), .B(n319), .X(n532));
sg13g2_a21oi_2 U1130 (.A1(net24685), .A2(N740), .B1(n1677), .Y(n1676));
sg13g2_nor2_2 U1131 (.A(n1678), .B(n4278), .Y(n1677));
sg13g2_a21oi_2 U1132 (.A1(net24743), .A2(N996), .B1(n1679), .Y(n1675));
sg13g2_nor2_2 U1133 (.A(n154), .B(n4282), .Y(n1679));
sg13g2_or2_1 U1134 (.A(n4281), .B(n318), .X(n531));
sg13g2_a21oi_2 U1135 (.A1(net24685), .A2(N741), .B1(n1682), .Y(n1681));
sg13g2_nor2_2 U1136 (.A(n1683), .B(n4278), .Y(n1682));
sg13g2_a21oi_2 U1137 (.A1(net24743), .A2(N997), .B1(n1684), .Y(n1680));
sg13g2_nor2_2 U1138 (.A(n153), .B(n4282), .Y(n1684));
sg13g2_or2_1 U1139 (.A(n4281), .B(n317), .X(n530));
sg13g2_a21oi_2 U1140 (.A1(n1134), .A2(N742), .B1(n1687), .Y(n1686));
sg13g2_nor2_2 U1141 (.A(n1688), .B(n4278), .Y(n1687));
sg13g2_a21oi_2 U1142 (.A1(net24743), .A2(N998), .B1(n1689), .Y(n1685));
sg13g2_nor2_2 U1143 (.A(n152), .B(n4282), .Y(n1689));
sg13g2_or2_1 U1144 (.A(n4281), .B(n298), .X(n529));
sg13g2_a21oi_2 U1145 (.A1(net24689), .A2(N743), .B1(n1692), .Y(n1691));
sg13g2_nor2_2 U1146 (.A(n1693), .B(n4278), .Y(n1692));
sg13g2_a21oi_2 U1147 (.A1(net24743), .A2(N999), .B1(n1694), .Y(n1690));
sg13g2_nor2_2 U1148 (.A(n151), .B(n4282), .Y(n1694));
sg13g2_or2_1 U1149 (.A(n4281), .B(n316), .X(n436));
sg13g2_a21oi_2 U1150 (.A1(net24687), .A2(N744), .B1(n1697), .Y(n1696));
sg13g2_nor2_2 U1151 (.A(n1698), .B(n4278), .Y(n1697));
sg13g2_a21oi_2 U1152 (.A1(net24743), .A2(N1000), .B1(n1699), .Y(n1695));
sg13g2_nor2_2 U1153 (.A(n150), .B(n4282), .Y(n1699));
sg13g2_or2_1 U1154 (.A(n4281), .B(n315), .X(n435));
sg13g2_a21oi_2 U1155 (.A1(net24685), .A2(N745), .B1(n1702), .Y(n1701));
sg13g2_nor2_2 U1156 (.A(n1703), .B(n4278), .Y(n1702));
sg13g2_a21oi_2 U1157 (.A1(net24743), .A2(N1001), .B1(n1704), .Y(n1700));
sg13g2_nor2_2 U1158 (.A(n149), .B(n4282), .Y(n1704));
sg13g2_or2_1 U1159 (.A(n4281), .B(n314), .X(n167));
sg13g2_a21oi_2 U1160 (.A1(net24687), .A2(N746), .B1(n1707), .Y(n1706));
sg13g2_nor2_2 U1161 (.A(n1708), .B(n4278), .Y(n1707));
sg13g2_a21oi_2 U1162 (.A1(net24743), .A2(N1002), .B1(n1709), .Y(n1705));
sg13g2_nor2_2 U1163 (.A(n148), .B(n4282), .Y(n1709));
sg13g2_or2_1 U1164 (.A(n4281), .B(n313), .X(n165));
sg13g2_a21oi_2 U1165 (.A1(net24689), .A2(N747), .B1(n1712), .Y(n1711));
sg13g2_nor2_2 U1166 (.A(n1713), .B(n4278), .Y(n1712));
sg13g2_a21oi_2 U1167 (.A1(net24743), .A2(N1003), .B1(n1714), .Y(n1710));
sg13g2_nor2_2 U1168 (.A(n147), .B(n4282), .Y(n1714));
sg13g2_or2_1 U1169 (.A(n4281), .B(n312), .X(n36));
sg13g2_a21oi_2 U1170 (.A1(net24687), .A2(N847), .B1(n1717), .Y(n1716));
sg13g2_nor2_2 U1171 (.A(n1718), .B(n4278), .Y(n1717));
sg13g2_a21oi_2 U1172 (.A1(net24743), .A2(N1103), .B1(n1719), .Y(n1715));
sg13g2_nor2_2 U1173 (.A(n47), .B(n4282), .Y(n1719));
sg13g2_or2_1 U1174 (.A(n4281), .B(n311), .X(n35));
sg13g2_a21oi_2 U1175 (.A1(net24689), .A2(N748), .B1(n1722), .Y(n1721));
sg13g2_nor2_2 U1176 (.A(n1723), .B(n4278), .Y(n1722));
sg13g2_a21oi_2 U1177 (.A1(net24743), .A2(N1004), .B1(n1724), .Y(n1720));
sg13g2_nor2_2 U1178 (.A(n146), .B(n4282), .Y(n1724));
sg13g2_or2_1 U1179 (.A(n4281), .B(n310), .X(n34));
sg13g2_a21oi_2 U1180 (.A1(n1134), .A2(N749), .B1(n1727), .Y(n1726));
sg13g2_nor2_2 U1181 (.A(n1728), .B(n4278), .Y(n1727));
sg13g2_a21oi_2 U1182 (.A1(net24743), .A2(N1005), .B1(n1729), .Y(n1725));
sg13g2_nor2_2 U1183 (.A(n145), .B(n4282), .Y(n1729));
sg13g2_or2_1 U1184 (.A(n4281), .B(n309), .X(n33));
sg13g2_a21oi_2 U1185 (.A1(net24685), .A2(N750), .B1(n1732), .Y(n1731));
sg13g2_nor2_2 U1186 (.A(n1733), .B(n4278), .Y(n1732));
sg13g2_a21oi_2 U1187 (.A1(net24743), .A2(N1006), .B1(n1734), .Y(n1730));
sg13g2_nor2_2 U1188 (.A(n144), .B(n4282), .Y(n1734));
sg13g2_or2_1 U1189 (.A(n4281), .B(n424), .X(n32));
sg13g2_a21oi_2 U1190 (.A1(net24685), .A2(N751), .B1(n1737), .Y(n1736));
sg13g2_nor2_2 U1191 (.A(n1738), .B(n4278), .Y(n1737));
sg13g2_a21oi_2 U1192 (.A1(net24743), .A2(N1007), .B1(n1739), .Y(n1735));
sg13g2_nor2_2 U1193 (.A(n143), .B(n4282), .Y(n1739));
sg13g2_or2_1 U1194 (.A(n4281), .B(n423), .X(n31));
sg13g2_a21oi_2 U1195 (.A1(net24689), .A2(N752), .B1(n1742), .Y(n1741));
sg13g2_nor2_2 U1196 (.A(n1743), .B(n4278), .Y(n1742));
sg13g2_a21oi_2 U1197 (.A1(net24743), .A2(N1008), .B1(n1744), .Y(n1740));
sg13g2_nor2_2 U1198 (.A(n142), .B(n4282), .Y(n1744));
sg13g2_or2_1 U1199 (.A(n4281), .B(n422), .X(n30));
sg13g2_a21oi_2 U1200 (.A1(net24685), .A2(N753), .B1(n1747), .Y(n1746));
sg13g2_nor2_2 U1201 (.A(n1748), .B(n4278), .Y(n1747));
sg13g2_a21oi_2 U1202 (.A1(net24743), .A2(N1009), .B1(n1749), .Y(n1745));
sg13g2_nor2_2 U1203 (.A(n141), .B(n4282), .Y(n1749));
sg13g2_or2_1 U1204 (.A(n4281), .B(n421), .X(n29));
sg13g2_a21oi_2 U1205 (.A1(net24687), .A2(N754), .B1(n1752), .Y(n1751));
sg13g2_nor2_2 U1206 (.A(n1753), .B(n4278), .Y(n1752));
sg13g2_a21oi_2 U1207 (.A1(net24743), .A2(N1010), .B1(n1754), .Y(n1750));
sg13g2_nor2_2 U1208 (.A(n140), .B(n4282), .Y(n1754));
sg13g2_or2_1 U1209 (.A(n4281), .B(n420), .X(n28));
sg13g2_a21oi_2 U1210 (.A1(net24685), .A2(N755), .B1(n1757), .Y(n1756));
sg13g2_nor2_2 U1211 (.A(n1758), .B(n4278), .Y(n1757));
sg13g2_a21oi_2 U1212 (.A1(net24743), .A2(N1011), .B1(n1759), .Y(n1755));
sg13g2_nor2_2 U1213 (.A(n139), .B(n4282), .Y(n1759));
sg13g2_or2_1 U1214 (.A(n4281), .B(n419), .X(n27));
sg13g2_a21oi_2 U1215 (.A1(net24687), .A2(N756), .B1(n1762), .Y(n1761));
sg13g2_nor2_2 U1216 (.A(n1763), .B(n4278), .Y(n1762));
sg13g2_a21oi_2 U1217 (.A1(net24743), .A2(N1012), .B1(n1764), .Y(n1760));
sg13g2_nor2_2 U1218 (.A(n138), .B(n4282), .Y(n1764));
sg13g2_or2_1 U1219 (.A(n4281), .B(n418), .X(n26));
sg13g2_a21oi_2 U1220 (.A1(net24685), .A2(N757), .B1(n1767), .Y(n1766));
sg13g2_nor2_2 U1221 (.A(n1768), .B(n4278), .Y(n1767));
sg13g2_a21oi_2 U1222 (.A1(net24743), .A2(N1013), .B1(n1769), .Y(n1765));
sg13g2_nor2_2 U1223 (.A(n137), .B(n4282), .Y(n1769));
sg13g2_or2_1 U1224 (.A(n4281), .B(n417), .X(n25));
sg13g2_a21oi_2 U1225 (.A1(net24685), .A2(N857), .B1(n1772), .Y(n1771));
sg13g2_nor2_2 U1226 (.A(n1773), .B(n4278), .Y(n1772));
sg13g2_a21oi_2 U1227 (.A1(net24743), .A2(N1113), .B1(n1774), .Y(n1770));
sg13g2_nor2_2 U1228 (.A(n37), .B(n4282), .Y(n1774));
sg13g2_or2_1 U1229 (.A(n4281), .B(n308), .X(n24));
sg13g2_or2_1 U1230 (.A(n4281), .B(n416), .X(n23));
sg13g2_or2_1 U1231 (.A(n4281), .B(n415), .X(n22));
sg13g2_o21ai_1 U1232 (.A1(n4327), .A2(n1136), .B1(n1776), .Y(mixcol_data_i_9));
sg13g2_nand2_2 U1233 (.A(subbytes_data_o_9), .B(n4317), .Y(n1776));
sg13g2_or2_1 U1234 (.A(n4281), .B(n414), .X(n21));
sg13g2_o21ai_1 U1235 (.A1(n4325), .A2(n1143), .B1(n1777), .Y(mixcol_data_i_99));
sg13g2_nand2_2 U1236 (.A(subbytes_data_o_99), .B(n4318), .Y(n1777));
sg13g2_or2_1 U1237 (.A(n4281), .B(n413), .X(n20));
sg13g2_o21ai_1 U1238 (.A1(n4328), .A2(n1148), .B1(n1778), .Y(mixcol_data_i_98));
sg13g2_nand2_2 U1239 (.A(subbytes_data_o_98), .B(n4321), .Y(n1778));
sg13g2_or2_1 U1240 (.A(n4281), .B(n412), .X(n19));
sg13g2_o21ai_1 U1241 (.A1(n4330), .A2(n1153), .B1(n1779), .Y(mixcol_data_i_97));
sg13g2_nand2_2 U1242 (.A(subbytes_data_o_97), .B(n4317), .Y(n1779));
sg13g2_or2_1 U1243 (.A(n4281), .B(n411), .X(n18));
sg13g2_o21ai_1 U1244 (.A1(n4328), .A2(n1158), .B1(n1780), .Y(mixcol_data_i_96));
sg13g2_nand2_2 U1245 (.A(subbytes_data_o_96), .B(n4321), .Y(n1780));
sg13g2_or2_1 U1246 (.A(n4281), .B(n410), .X(n17));
sg13g2_o21ai_1 U1247 (.A1(n4328), .A2(n1163), .B1(n1781), .Y(mixcol_data_i_95));
sg13g2_nand2_2 U1248 (.A(subbytes_data_o_95), .B(n4316), .Y(n1781));
sg13g2_or2_1 U1249 (.A(n4281), .B(n409), .X(n16));
sg13g2_o21ai_1 U1250 (.A1(n4328), .A2(n1168), .B1(n1782), .Y(mixcol_data_i_94));
sg13g2_nand2_2 U1251 (.A(subbytes_data_o_94), .B(n4318), .Y(n1782));
sg13g2_or2_1 U1252 (.A(n4281), .B(n408), .X(n15));
sg13g2_o21ai_1 U1253 (.A1(n4328), .A2(n1173), .B1(n1783), .Y(mixcol_data_i_93));
sg13g2_nand2_2 U1254 (.A(subbytes_data_o_93), .B(n4318), .Y(n1783));
sg13g2_or2_1 U1255 (.A(n4281), .B(n407), .X(n14));
sg13g2_o21ai_1 U1256 (.A1(n4328), .A2(n1178), .B1(n1784), .Y(mixcol_data_i_92));
sg13g2_nand2_2 U1257 (.A(subbytes_data_o_92), .B(n4316), .Y(n1784));
sg13g2_or2_1 U1258 (.A(n4281), .B(n307), .X(n13));
sg13g2_o21ai_1 U1259 (.A1(n4328), .A2(n1183), .B1(n1785), .Y(mixcol_data_i_91));
sg13g2_nand2_2 U1260 (.A(subbytes_data_o_91), .B(n4316), .Y(n1785));
sg13g2_or2_1 U1261 (.A(n4281), .B(n406), .X(n12));
sg13g2_o21ai_1 U1262 (.A1(n4328), .A2(n1188), .B1(n1786), .Y(mixcol_data_i_90));
sg13g2_nand2_2 U1263 (.A(subbytes_data_o_90), .B(n4319), .Y(n1786));
sg13g2_or2_1 U1264 (.A(n4281), .B(n405), .X(n11));
sg13g2_o21ai_1 U1265 (.A1(n4328), .A2(n1193), .B1(n1787), .Y(mixcol_data_i_8));
sg13g2_nand2_2 U1266 (.A(subbytes_data_o_8), .B(n4316), .Y(n1787));
sg13g2_or2_1 U1267 (.A(n4281), .B(n404), .X(n10));
sg13g2_o21ai_1 U1268 (.A1(n4328), .A2(n1198), .B1(n1788), .Y(mixcol_data_i_89));
sg13g2_nand2_2 U1269 (.A(subbytes_data_o_89), .B(n4318), .Y(n1788));
sg13g2_or2_1 U1270 (.A(n4281), .B(n403), .X(n9));
sg13g2_o21ai_1 U1271 (.A1(n4328), .A2(n1203), .B1(n1789), .Y(mixcol_data_i_88));
sg13g2_nand2_2 U1272 (.A(subbytes_data_o_88), .B(n4318), .Y(n1789));
sg13g2_or2_1 U1273 (.A(n4281), .B(n402), .X(n8));
sg13g2_o21ai_1 U1274 (.A1(n4328), .A2(n1208), .B1(n1790), .Y(mixcol_data_i_87));
sg13g2_nand2_2 U1275 (.A(subbytes_data_o_87), .B(n4319), .Y(n1790));
sg13g2_or2_1 U1276 (.A(n4281), .B(n401), .X(n7));
sg13g2_o21ai_1 U1277 (.A1(n4329), .A2(n1213), .B1(n1791), .Y(mixcol_data_i_86));
sg13g2_nand2_2 U1278 (.A(subbytes_data_o_86), .B(n4317), .Y(n1791));
sg13g2_or2_1 U1279 (.A(n4281), .B(n400), .X(n6));
sg13g2_o21ai_1 U1280 (.A1(n4329), .A2(n1218), .B1(n1792), .Y(mixcol_data_i_85));
sg13g2_nand2_2 U1281 (.A(subbytes_data_o_85), .B(n4318), .Y(n1792));
sg13g2_or2_1 U1282 (.A(n4281), .B(n399), .X(n5));
sg13g2_o21ai_1 U1283 (.A1(n4326), .A2(n1223), .B1(n1793), .Y(mixcol_data_i_84));
sg13g2_nand2_2 U1284 (.A(subbytes_data_o_84), .B(n4319), .Y(n1793));
sg13g2_or2_1 U1285 (.A(n4281), .B(n398), .X(n4));
sg13g2_o21ai_1 U1286 (.A1(n4325), .A2(n1228), .B1(n1794), .Y(mixcol_data_i_83));
sg13g2_nand2_2 U1287 (.A(subbytes_data_o_83), .B(n4319), .Y(n1794));
sg13g2_or2_1 U1288 (.A(n4281), .B(n397), .X(n3));
sg13g2_o21ai_1 U1289 (.A1(n4327), .A2(n1233), .B1(n1795), .Y(mixcol_data_i_82));
sg13g2_nand2_2 U1290 (.A(subbytes_data_o_82), .B(n4320), .Y(n1795));
sg13g2_or2_1 U1291 (.A(n4281), .B(n297), .X(n2));
sg13g2_o21ai_1 U1292 (.A1(n4328), .A2(n1238), .B1(n1796), .Y(mixcol_data_i_81));
sg13g2_nand2_2 U1293 (.A(subbytes_data_o_81), .B(n4318), .Y(n1796));
sg13g2_o21ai_1 U1295 (.A1(n4329), .A2(n1243), .B1(n1797), .Y(mixcol_data_i_80));
sg13g2_nand2_2 U1296 (.A(subbytes_data_o_80), .B(n4317), .Y(n1797));
sg13g2_o21ai_1 U1298 (.A1(n4326), .A2(n1248), .B1(n1798), .Y(mixcol_data_i_7));
sg13g2_nand2_2 U1299 (.A(subbytes_data_o_7), .B(n4318), .Y(n1798));
sg13g2_o21ai_1 U1301 (.A1(n4326), .A2(n1253), .B1(n1799), .Y(mixcol_data_i_79));
sg13g2_nand2_2 U1302 (.A(subbytes_data_o_79), .B(n4318), .Y(n1799));
sg13g2_o21ai_1 U1304 (.A1(n4328), .A2(n1258), .B1(n1800), .Y(mixcol_data_i_78));
sg13g2_nand2_2 U1305 (.A(subbytes_data_o_78), .B(n4317), .Y(n1800));
sg13g2_o21ai_1 U1307 (.A1(n4325), .A2(n1263), .B1(n1801), .Y(mixcol_data_i_77));
sg13g2_nand2_2 U1308 (.A(subbytes_data_o_77), .B(n4317), .Y(n1801));
sg13g2_o21ai_1 U1310 (.A1(n4329), .A2(n1268), .B1(n1802), .Y(mixcol_data_i_76));
sg13g2_nand2_2 U1311 (.A(subbytes_data_o_76), .B(n4318), .Y(n1802));
sg13g2_o21ai_1 U1313 (.A1(n4329), .A2(n1273), .B1(n1803), .Y(mixcol_data_i_75));
sg13g2_nand2_2 U1314 (.A(subbytes_data_o_75), .B(n4318), .Y(n1803));
sg13g2_o21ai_1 U1316 (.A1(n4329), .A2(n1278), .B1(n1804), .Y(mixcol_data_i_74));
sg13g2_nand2_2 U1317 (.A(subbytes_data_o_74), .B(n4316), .Y(n1804));
sg13g2_o21ai_1 U1319 (.A1(n4329), .A2(n1283), .B1(n1805), .Y(mixcol_data_i_73));
sg13g2_nand2_2 U1320 (.A(subbytes_data_o_73), .B(n4319), .Y(n1805));
sg13g2_o21ai_1 U1322 (.A1(n4329), .A2(n1288), .B1(n1806), .Y(mixcol_data_i_72));
sg13g2_nand2_2 U1323 (.A(subbytes_data_o_72), .B(n4298), .Y(n1806));
sg13g2_o21ai_1 U1325 (.A1(n4329), .A2(n1293), .B1(n1807), .Y(mixcol_data_i_71));
sg13g2_nand2_2 U1326 (.A(subbytes_data_o_71), .B(n4323), .Y(n1807));
sg13g2_o21ai_1 U1328 (.A1(n4329), .A2(n1298), .B1(n1808), .Y(mixcol_data_i_70));
sg13g2_nand2_2 U1329 (.A(subbytes_data_o_70), .B(n4298), .Y(n1808));
sg13g2_o21ai_1 U1331 (.A1(n4329), .A2(n1303), .B1(n1809), .Y(mixcol_data_i_6));
sg13g2_nand2_2 U1332 (.A(subbytes_data_o_6), .B(n4318), .Y(n1809));
sg13g2_o21ai_1 U1334 (.A1(n4329), .A2(n1308), .B1(n1810), .Y(mixcol_data_i_69));
sg13g2_nand2_2 U1335 (.A(subbytes_data_o_69), .B(n4317), .Y(n1810));
sg13g2_o21ai_1 U1337 (.A1(n4329), .A2(n1313), .B1(n1811), .Y(mixcol_data_i_68));
sg13g2_nand2_2 U1338 (.A(subbytes_data_o_68), .B(n4298), .Y(n1811));
sg13g2_o21ai_1 U1340 (.A1(n4329), .A2(n1318), .B1(n1812), .Y(mixcol_data_i_67));
sg13g2_nand2_2 U1341 (.A(subbytes_data_o_67), .B(n4316), .Y(n1812));
sg13g2_o21ai_1 U1343 (.A1(n4327), .A2(n1323), .B1(n1813), .Y(mixcol_data_i_66));
sg13g2_nand2_2 U1344 (.A(subbytes_data_o_66), .B(n4318), .Y(n1813));
sg13g2_o21ai_1 U1346 (.A1(n4328), .A2(n1328), .B1(n1814), .Y(mixcol_data_i_65));
sg13g2_nand2_2 U1347 (.A(subbytes_data_o_65), .B(n4318), .Y(n1814));
sg13g2_o21ai_1 U1349 (.A1(n4327), .A2(n1333), .B1(n1815), .Y(mixcol_data_i_64));
sg13g2_nand2_2 U1350 (.A(subbytes_data_o_64), .B(n4321), .Y(n1815));
sg13g2_nand2_2 U1353 (.A(subbytes_data_o_63), .B(n4321), .Y(n1816));
sg13g2_o21ai_1 U1355 (.A1(n4328), .A2(n1343), .B1(n1817), .Y(mixcol_data_i_62));
sg13g2_nand2_2 U1356 (.A(subbytes_data_o_62), .B(n4298), .Y(n1817));
sg13g2_o21ai_1 U1358 (.A1(n4325), .A2(n1348), .B1(n1818), .Y(mixcol_data_i_61));
sg13g2_o21ai_1 U1361 (.A1(n4329), .A2(n1353), .B1(n1819), .Y(mixcol_data_i_60));
sg13g2_nand2_2 U1362 (.A(subbytes_data_o_60), .B(n4318), .Y(n1819));
sg13g2_o21ai_1 U1364 (.A1(n4328), .A2(n1358), .B1(n1820), .Y(mixcol_data_i_5));
sg13g2_nand2_2 U1365 (.A(subbytes_data_o_5), .B(n4320), .Y(n1820));
sg13g2_o21ai_1 U1367 (.A1(n4326), .A2(n1363), .B1(n1821), .Y(mixcol_data_i_59));
sg13g2_nand2_2 U1368 (.A(subbytes_data_o_59), .B(n4319), .Y(n1821));
sg13g2_o21ai_1 U1370 (.A1(n4326), .A2(n1368), .B1(n1822), .Y(mixcol_data_i_58));
sg13g2_nand2_2 U1371 (.A(subbytes_data_o_58), .B(n4321), .Y(n1822));
sg13g2_o21ai_1 U1373 (.A1(n4330), .A2(n1373), .B1(n1823), .Y(mixcol_data_i_57));
sg13g2_nand2_2 U1374 (.A(subbytes_data_o_57), .B(n4321), .Y(n1823));
sg13g2_o21ai_1 U1376 (.A1(n4330), .A2(n1378), .B1(n1824), .Y(mixcol_data_i_56));
sg13g2_nand2_2 U1377 (.A(subbytes_data_o_56), .B(n4317), .Y(n1824));
sg13g2_o21ai_1 U1379 (.A1(n4330), .A2(n1383), .B1(n1825), .Y(mixcol_data_i_55));
sg13g2_o21ai_1 U1382 (.A1(n4330), .A2(n1388), .B1(n1826), .Y(mixcol_data_i_54));
sg13g2_nand2_2 U1383 (.A(subbytes_data_o_54), .B(n4319), .Y(n1826));
sg13g2_o21ai_1 U1385 (.A1(n4330), .A2(n1393), .B1(n1827), .Y(mixcol_data_i_53));
sg13g2_o21ai_1 U1388 (.A1(n4330), .A2(n1398), .B1(n1828), .Y(mixcol_data_i_52));
sg13g2_nand2_2 U1389 (.A(subbytes_data_o_52), .B(n4320), .Y(n1828));
sg13g2_o21ai_1 U1391 (.A1(n4330), .A2(n1403), .B1(n1829), .Y(mixcol_data_i_51));
sg13g2_o21ai_1 U1394 (.A1(n4330), .A2(n1408), .B1(n1830), .Y(mixcol_data_i_50));
sg13g2_nand2_2 U1395 (.A(subbytes_data_o_50), .B(n4320), .Y(n1830));
sg13g2_o21ai_1 U1397 (.A1(n4330), .A2(n1413), .B1(n1831), .Y(mixcol_data_i_4));
sg13g2_nand2_2 U1398 (.A(subbytes_data_o_4), .B(n4320), .Y(n1831));
sg13g2_o21ai_1 U1400 (.A1(n4330), .A2(n1418), .B1(n1832), .Y(mixcol_data_i_49));
sg13g2_o21ai_1 U1403 (.A1(n4330), .A2(n1423), .B1(n1833), .Y(mixcol_data_i_48));
sg13g2_nand2_2 U1404 (.A(subbytes_data_o_48), .B(n4320), .Y(n1833));
sg13g2_o21ai_1 U1406 (.A1(n4330), .A2(n1428), .B1(n1834), .Y(mixcol_data_i_47));
sg13g2_o21ai_1 U1409 (.A1(n4329), .A2(n1433), .B1(n1835), .Y(mixcol_data_i_46));
sg13g2_o21ai_1 U1412 (.A1(n4327), .A2(n1438), .B1(n1836), .Y(mixcol_data_i_45));
sg13g2_nand2_2 U1413 (.A(subbytes_data_o_45), .B(n4320), .Y(n1836));
sg13g2_o21ai_1 U1415 (.A1(n4326), .A2(n1443), .B1(n1837), .Y(mixcol_data_i_44));
sg13g2_nand2_2 U1416 (.A(subbytes_data_o_44), .B(n4320), .Y(n1837));
sg13g2_o21ai_1 U1418 (.A1(n4325), .A2(n1448), .B1(n1838), .Y(mixcol_data_i_43));
sg13g2_nand2_2 U1419 (.A(subbytes_data_o_43), .B(n4319), .Y(n1838));
sg13g2_o21ai_1 U1421 (.A1(n4327), .A2(n1453), .B1(n1839), .Y(mixcol_data_i_42));
sg13g2_nand2_2 U1422 (.A(subbytes_data_o_42), .B(n4319), .Y(n1839));
sg13g2_o21ai_1 U1424 (.A1(n4328), .A2(n1458), .B1(n1840), .Y(mixcol_data_i_41));
sg13g2_nand2_2 U1425 (.A(subbytes_data_o_41), .B(n4319), .Y(n1840));
sg13g2_o21ai_1 U1427 (.A1(n4330), .A2(n1463), .B1(n1841), .Y(mixcol_data_i_40));
sg13g2_o21ai_1 U1430 (.A1(n4325), .A2(n1468), .B1(n1842), .Y(mixcol_data_i_3));
sg13g2_nand2_2 U1431 (.A(subbytes_data_o_3), .B(n4319), .Y(n1842));
sg13g2_o21ai_1 U1433 (.A1(n4328), .A2(n1473), .B1(n1843), .Y(mixcol_data_i_39));
sg13g2_nand2_2 U1434 (.A(subbytes_data_o_39), .B(n4319), .Y(n1843));
sg13g2_o21ai_1 U1436 (.A1(n4327), .A2(n1478), .B1(n1844), .Y(mixcol_data_i_38));
sg13g2_nand2_2 U1437 (.A(subbytes_data_o_38), .B(n4319), .Y(n1844));
sg13g2_o21ai_1 U1439 (.A1(n4328), .A2(n1483), .B1(n1845), .Y(mixcol_data_i_37));
sg13g2_nand2_2 U1440 (.A(subbytes_data_o_37), .B(n4319), .Y(n1845));
sg13g2_o21ai_1 U1442 (.A1(n4326), .A2(n1488), .B1(n1846), .Y(mixcol_data_i_36));
sg13g2_nand2_2 U1443 (.A(subbytes_data_o_36), .B(n4319), .Y(n1846));
sg13g2_o21ai_1 U1445 (.A1(n4326), .A2(n1493), .B1(n1847), .Y(mixcol_data_i_35));
sg13g2_nand2_2 U1446 (.A(subbytes_data_o_35), .B(n4319), .Y(n1847));
sg13g2_o21ai_1 U1448 (.A1(n4328), .A2(n1498), .B1(n1848), .Y(mixcol_data_i_34));
sg13g2_nand2_2 U1449 (.A(subbytes_data_o_34), .B(n4319), .Y(n1848));
sg13g2_o21ai_1 U1451 (.A1(n4329), .A2(n1503), .B1(n1849), .Y(mixcol_data_i_33));
sg13g2_nand2_2 U1452 (.A(subbytes_data_o_33), .B(n4318), .Y(n1849));
sg13g2_o21ai_1 U1454 (.A1(n4330), .A2(n1508), .B1(n1850), .Y(mixcol_data_i_32));
sg13g2_nand2_2 U1455 (.A(subbytes_data_o_32), .B(n4298), .Y(n1850));
sg13g2_o21ai_1 U1457 (.A1(n4327), .A2(n1513), .B1(n1851), .Y(mixcol_data_i_31));
sg13g2_nand2_2 U1458 (.A(subbytes_data_o_31), .B(n4321), .Y(n1851));
sg13g2_o21ai_1 U1460 (.A1(n4326), .A2(n1518), .B1(n1852), .Y(mixcol_data_i_30));
sg13g2_nand2_2 U1461 (.A(subbytes_data_o_30), .B(n4318), .Y(n1852));
sg13g2_o21ai_1 U1463 (.A1(n4330), .A2(n1523), .B1(n1853), .Y(mixcol_data_i_2));
sg13g2_nand2_2 U1464 (.A(subbytes_data_o_2), .B(n4321), .Y(n1853));
sg13g2_o21ai_1 U1466 (.A1(n4327), .A2(n1528), .B1(n1854), .Y(mixcol_data_i_29));
sg13g2_o21ai_1 U1469 (.A1(n4330), .A2(n1533), .B1(n1855), .Y(mixcol_data_i_28));
sg13g2_nand2_2 U1470 (.A(subbytes_data_o_28), .B(n4321), .Y(n1855));
sg13g2_o21ai_1 U1472 (.A1(n4328), .A2(n1538), .B1(n1856), .Y(mixcol_data_i_27));
sg13g2_nand2_2 U1473 (.A(subbytes_data_o_27), .B(n4298), .Y(n1856));
sg13g2_o21ai_1 U1475 (.A1(n4329), .A2(n1543), .B1(n1857), .Y(mixcol_data_i_26));
sg13g2_nand2_2 U1476 (.A(subbytes_data_o_26), .B(n4317), .Y(n1857));
sg13g2_o21ai_1 U1478 (.A1(n4329), .A2(n1548), .B1(n1858), .Y(mixcol_data_i_25));
sg13g2_nand2_2 U1479 (.A(subbytes_data_o_25), .B(n4298), .Y(n1858));
sg13g2_o21ai_1 U1481 (.A1(n4329), .A2(n1553), .B1(n1859), .Y(mixcol_data_i_24));
sg13g2_nand2_2 U1482 (.A(subbytes_data_o_24), .B(n4319), .Y(n1859));
sg13g2_o21ai_1 U1484 (.A1(n4326), .A2(n1558), .B1(n1860), .Y(mixcol_data_i_23));
sg13g2_nand2_2 U1485 (.A(subbytes_data_o_23), .B(n4318), .Y(n1860));
sg13g2_o21ai_1 U1487 (.A1(n4329), .A2(n1563), .B1(n1861), .Y(mixcol_data_i_22));
sg13g2_nand2_2 U1488 (.A(subbytes_data_o_22), .B(n4318), .Y(n1861));
sg13g2_o21ai_1 U1490 (.A1(n4326), .A2(n1568), .B1(n1862), .Y(mixcol_data_i_21));
sg13g2_o21ai_1 U1493 (.A1(n4328), .A2(n1573), .B1(n1863), .Y(mixcol_data_i_20));
sg13g2_nand2_2 U1494 (.A(subbytes_data_o_20), .B(n4318), .Y(n1863));
sg13g2_o21ai_1 U1496 (.A1(n4326), .A2(n1578), .B1(n1864), .Y(mixcol_data_i_1));
sg13g2_nand2_2 U1497 (.A(subbytes_data_o_1), .B(n4318), .Y(n1864));
sg13g2_o21ai_1 U1499 (.A1(n4328), .A2(n1583), .B1(n1865), .Y(mixcol_data_i_19));
sg13g2_nand2_2 U1500 (.A(subbytes_data_o_19), .B(n4318), .Y(n1865));
sg13g2_o21ai_1 U1502 (.A1(n4330), .A2(n1588), .B1(n1866), .Y(mixcol_data_i_18));
sg13g2_nand2_2 U1503 (.A(subbytes_data_o_18), .B(n4318), .Y(n1866));
sg13g2_o21ai_1 U1505 (.A1(n4330), .A2(n1593), .B1(n1867), .Y(mixcol_data_i_17));
sg13g2_nand2_2 U1506 (.A(subbytes_data_o_17), .B(n4318), .Y(n1867));
sg13g2_o21ai_1 U1508 (.A1(n4330), .A2(n1598), .B1(n1868), .Y(mixcol_data_i_16));
sg13g2_nand2_2 U1509 (.A(subbytes_data_o_16), .B(n4318), .Y(n1868));
sg13g2_o21ai_1 U1511 (.A1(n4330), .A2(n1603), .B1(n1869), .Y(mixcol_data_i_15));
sg13g2_nand2_2 U1512 (.A(subbytes_data_o_15), .B(n4318), .Y(n1869));
sg13g2_o21ai_1 U1514 (.A1(n4328), .A2(n1608), .B1(n1870), .Y(mixcol_data_i_14));
sg13g2_nand2_2 U1515 (.A(subbytes_data_o_14), .B(n4318), .Y(n1870));
sg13g2_o21ai_1 U1517 (.A1(n4329), .A2(n1613), .B1(n1871), .Y(mixcol_data_i_13));
sg13g2_nand2_2 U1518 (.A(subbytes_data_o_13), .B(n4317), .Y(n1871));
sg13g2_o21ai_1 U1520 (.A1(n4325), .A2(n1618), .B1(n1872), .Y(mixcol_data_i_12));
sg13g2_nand2_2 U1521 (.A(subbytes_data_o_12), .B(n4318), .Y(n1872));
sg13g2_o21ai_1 U1523 (.A1(n4330), .A2(n1623), .B1(n1873), .Y(mixcol_data_i_127));
sg13g2_nand2_2 U1524 (.A(subbytes_data_o_127), .B(n4318), .Y(n1873));
sg13g2_o21ai_1 U1526 (.A1(n4328), .A2(n1628), .B1(n1874), .Y(mixcol_data_i_126));
sg13g2_nand2_2 U1527 (.A(subbytes_data_o_126), .B(n4317), .Y(n1874));
sg13g2_o21ai_1 U1529 (.A1(n4328), .A2(n1633), .B1(n1875), .Y(mixcol_data_i_125));
sg13g2_nand2_2 U1530 (.A(subbytes_data_o_125), .B(n4318), .Y(n1875));
sg13g2_o21ai_1 U1532 (.A1(n4330), .A2(n1638), .B1(n1876), .Y(mixcol_data_i_124));
sg13g2_nand2_2 U1533 (.A(subbytes_data_o_124), .B(n4316), .Y(n1876));
sg13g2_o21ai_1 U1535 (.A1(n4328), .A2(n1643), .B1(n1877), .Y(mixcol_data_i_123));
sg13g2_nand2_2 U1536 (.A(subbytes_data_o_123), .B(n4316), .Y(n1877));
sg13g2_o21ai_1 U1538 (.A1(n4329), .A2(n1648), .B1(n1878), .Y(mixcol_data_i_122));
sg13g2_nand2_2 U1539 (.A(subbytes_data_o_122), .B(n4317), .Y(n1878));
sg13g2_o21ai_1 U1541 (.A1(n4326), .A2(n1653), .B1(n1879), .Y(mixcol_data_i_121));
sg13g2_nand2_2 U1542 (.A(subbytes_data_o_121), .B(n4316), .Y(n1879));
sg13g2_o21ai_1 U1544 (.A1(n4327), .A2(n1658), .B1(n1880), .Y(mixcol_data_i_120));
sg13g2_nand2_2 U1545 (.A(subbytes_data_o_120), .B(n4318), .Y(n1880));
sg13g2_o21ai_1 U1547 (.A1(n4330), .A2(n1663), .B1(n1881), .Y(mixcol_data_i_11));
sg13g2_nand2_2 U1548 (.A(subbytes_data_o_11), .B(n4318), .Y(n1881));
sg13g2_o21ai_1 U1550 (.A1(n4328), .A2(n1668), .B1(n1882), .Y(mixcol_data_i_119));
sg13g2_nand2_2 U1551 (.A(subbytes_data_o_119), .B(n4317), .Y(n1882));
sg13g2_o21ai_1 U1553 (.A1(n4330), .A2(n1673), .B1(n1883), .Y(mixcol_data_i_118));
sg13g2_nand2_2 U1554 (.A(subbytes_data_o_118), .B(n4317), .Y(n1883));
sg13g2_o21ai_1 U1556 (.A1(n4325), .A2(n1678), .B1(n1884), .Y(mixcol_data_i_117));
sg13g2_nand2_2 U1557 (.A(subbytes_data_o_117), .B(n4317), .Y(n1884));
sg13g2_o21ai_1 U1559 (.A1(n4330), .A2(n1683), .B1(n1885), .Y(mixcol_data_i_116));
sg13g2_nand2_2 U1560 (.A(subbytes_data_o_116), .B(n4317), .Y(n1885));
sg13g2_o21ai_1 U1562 (.A1(n4328), .A2(n1688), .B1(n1886), .Y(mixcol_data_i_115));
sg13g2_nand2_2 U1563 (.A(subbytes_data_o_115), .B(n4317), .Y(n1886));
sg13g2_o21ai_1 U1565 (.A1(n4327), .A2(n1693), .B1(n1887), .Y(mixcol_data_i_114));
sg13g2_nand2_2 U1566 (.A(subbytes_data_o_114), .B(n4317), .Y(n1887));
sg13g2_o21ai_1 U1568 (.A1(n4329), .A2(n1698), .B1(n1888), .Y(mixcol_data_i_113));
sg13g2_nand2_2 U1569 (.A(subbytes_data_o_113), .B(n4317), .Y(n1888));
sg13g2_o21ai_1 U1571 (.A1(n4325), .A2(n1703), .B1(n1889), .Y(mixcol_data_i_112));
sg13g2_nand2_2 U1572 (.A(subbytes_data_o_112), .B(n4317), .Y(n1889));
sg13g2_o21ai_1 U1574 (.A1(n4326), .A2(n1708), .B1(n1890), .Y(mixcol_data_i_111));
sg13g2_nand2_2 U1575 (.A(subbytes_data_o_111), .B(n4317), .Y(n1890));
sg13g2_o21ai_1 U1577 (.A1(n4330), .A2(n1713), .B1(n1891), .Y(mixcol_data_i_110));
sg13g2_nand2_2 U1578 (.A(subbytes_data_o_110), .B(n4317), .Y(n1891));
sg13g2_o21ai_1 U1580 (.A1(n4330), .A2(n1718), .B1(n1892), .Y(mixcol_data_i_10));
sg13g2_nand2_2 U1581 (.A(subbytes_data_o_10), .B(n4317), .Y(n1892));
sg13g2_o21ai_1 U1583 (.A1(n4329), .A2(n1723), .B1(n1893), .Y(mixcol_data_i_109));
sg13g2_nand2_2 U1584 (.A(subbytes_data_o_109), .B(n4316), .Y(n1893));
sg13g2_o21ai_1 U1586 (.A1(n4330), .A2(n1728), .B1(n1894), .Y(mixcol_data_i_108));
sg13g2_nand2_2 U1587 (.A(subbytes_data_o_108), .B(n4316), .Y(n1894));
sg13g2_o21ai_1 U1589 (.A1(n4326), .A2(n1733), .B1(n1895), .Y(mixcol_data_i_107));
sg13g2_nand2_2 U1590 (.A(subbytes_data_o_107), .B(n4316), .Y(n1895));
sg13g2_o21ai_1 U1592 (.A1(n4329), .A2(n1738), .B1(n1896), .Y(mixcol_data_i_106));
sg13g2_nand2_2 U1593 (.A(subbytes_data_o_106), .B(n4316), .Y(n1896));
sg13g2_o21ai_1 U1595 (.A1(n4330), .A2(n1743), .B1(n1897), .Y(mixcol_data_i_105));
sg13g2_nand2_2 U1596 (.A(subbytes_data_o_105), .B(n4316), .Y(n1897));
sg13g2_o21ai_1 U1598 (.A1(n4327), .A2(n1748), .B1(n1898), .Y(mixcol_data_i_104));
sg13g2_nand2_2 U1599 (.A(subbytes_data_o_104), .B(n4316), .Y(n1898));
sg13g2_o21ai_1 U1601 (.A1(n4326), .A2(n1753), .B1(n1899), .Y(mixcol_data_i_103));
sg13g2_o21ai_1 U1604 (.A1(n4330), .A2(n1758), .B1(n1900), .Y(mixcol_data_i_102));
sg13g2_nand2_2 U1605 (.A(subbytes_data_o_102), .B(n4316), .Y(n1900));
sg13g2_o21ai_1 U1607 (.A1(n4327), .A2(n1763), .B1(n1901), .Y(mixcol_data_i_101));
sg13g2_nand2_2 U1608 (.A(subbytes_data_o_101), .B(n4316), .Y(n1901));
sg13g2_o21ai_1 U1610 (.A1(n4327), .A2(n1768), .B1(n1902), .Y(mixcol_data_i_100));
sg13g2_nand2_2 U1611 (.A(subbytes_data_o_100), .B(n4316), .Y(n1902));
sg13g2_o21ai_1 U1613 (.A1(n4326), .A2(n1773), .B1(n1903), .Y(mixcol_data_i_0));
sg13g2_nand2_2 U1614 (.A(subbytes_data_o_0), .B(n4316), .Y(n1903));
sg13g2_nand2_2 U1619 (.A(n4212), .B(N1538), .Y(n1907));
sg13g2_nand2_2 U1623 (.A(n4212), .B(N1536), .Y(n1910));
sg13g2_inv_4 U1629 (.A(key_i_9_), .Y(n852));
sg13g2_o21ai_1 U1630 (.A1(n4221), .A2(n1917), .B1(n1918), .Y(keysched_last_key_i_99));
sg13g2_nand2_2 U1631 (.A(keysched_new_key_o_99), .B(net25892), .Y(n1918));
sg13g2_inv_4 U1632 (.A(key_i_99_), .Y(n1917));
sg13g2_o21ai_1 U1633 (.A1(net26188), .A2(n1919), .B1(n1920), .Y(keysched_last_key_i_98));
sg13g2_nand2_2 U1634 (.A(keysched_new_key_o_98), .B(net25892), .Y(n1920));
sg13g2_inv_4 U1635 (.A(key_i_98_), .Y(n1919));
sg13g2_o21ai_1 U1636 (.A1(n4221), .A2(n1921), .B1(n1922), .Y(keysched_last_key_i_97));
sg13g2_nand2_2 U1637 (.A(keysched_new_key_o_97), .B(net25895), .Y(n1922));
sg13g2_inv_4 U1638 (.A(key_i_97_), .Y(n1921));
sg13g2_nand2_2 U1640 (.A(keysched_new_key_o_96), .B(net25895), .Y(n1924));
sg13g2_inv_4 U1641 (.A(key_i_96_), .Y(n1923));
sg13g2_o21ai_1 U1642 (.A1(n4221), .A2(n1925), .B1(n1926), .Y(keysched_last_key_i_95));
sg13g2_nand2_2 U1643 (.A(keysched_new_key_o_95), .B(n4155), .Y(n1926));
sg13g2_inv_4 U1644 (.A(key_i_95_), .Y(n1925));
sg13g2_o21ai_1 U1645 (.A1(n4221), .A2(n1927), .B1(n1928), .Y(keysched_last_key_i_94));
sg13g2_nand2_2 U1646 (.A(keysched_new_key_o_94), .B(n4155), .Y(n1928));
sg13g2_inv_4 U1647 (.A(key_i_94_), .Y(n1927));
sg13g2_o21ai_1 U1648 (.A1(net26188), .A2(n1929), .B1(n1930), .Y(keysched_last_key_i_93));
sg13g2_nand2_2 U1649 (.A(keysched_new_key_o_93), .B(n4155), .Y(n1930));
sg13g2_inv_4 U1650 (.A(key_i_93_), .Y(n1929));
sg13g2_o21ai_1 U1651 (.A1(n4221), .A2(n1931), .B1(n1932), .Y(keysched_last_key_i_92));
sg13g2_nand2_2 U1652 (.A(keysched_new_key_o_92), .B(net24851), .Y(n1932));
sg13g2_inv_4 U1653 (.A(key_i_92_), .Y(n1931));
sg13g2_o21ai_1 U1654 (.A1(net26188), .A2(n1933), .B1(n1934), .Y(keysched_last_key_i_91));
sg13g2_nand2_2 U1655 (.A(keysched_new_key_o_91), .B(net24851), .Y(n1934));
sg13g2_inv_4 U1656 (.A(key_i_91_), .Y(n1933));
sg13g2_o21ai_1 U1657 (.A1(n4221), .A2(n1935), .B1(n1936), .Y(keysched_last_key_i_90));
sg13g2_nand2_2 U1658 (.A(keysched_new_key_o_90), .B(net24847), .Y(n1936));
sg13g2_inv_4 U1659 (.A(key_i_90_), .Y(n1935));
sg13g2_inv_4 U1662 (.A(key_i_8_), .Y(n858));
sg13g2_nand2_2 U1664 (.A(keysched_new_key_o_89), .B(net26430), .Y(n1939));
sg13g2_inv_4 U1665 (.A(key_i_89_), .Y(n1938));
sg13g2_o21ai_1 U1666 (.A1(net26188), .A2(n1940), .B1(n1941), .Y(keysched_last_key_i_88));
sg13g2_nand2_2 U1667 (.A(keysched_new_key_o_88), .B(n4156), .Y(n1941));
sg13g2_inv_4 U1668 (.A(key_i_88_), .Y(n1940));
sg13g2_o21ai_1 U1669 (.A1(net24783), .A2(n1942), .B1(n1943), .Y(keysched_last_key_i_87));
sg13g2_nand2_2 U1670 (.A(keysched_new_key_o_87), .B(n4156), .Y(n1943));
sg13g2_inv_4 U1671 (.A(key_i_87_), .Y(n1942));
sg13g2_o21ai_1 U1672 (.A1(net26188), .A2(n1944), .B1(n1945), .Y(keysched_last_key_i_86));
sg13g2_nand2_2 U1673 (.A(keysched_new_key_o_86), .B(net25895), .Y(n1945));
sg13g2_inv_4 U1674 (.A(key_i_86_), .Y(n1944));
sg13g2_o21ai_1 U1675 (.A1(net24795), .A2(n1946), .B1(n1947), .Y(keysched_last_key_i_85));
sg13g2_nand2_2 U1676 (.A(keysched_new_key_o_85), .B(net24845), .Y(n1947));
sg13g2_inv_4 U1677 (.A(key_i_85_), .Y(n1946));
sg13g2_o21ai_1 U1678 (.A1(net26188), .A2(n1948), .B1(n1949), .Y(keysched_last_key_i_84));
sg13g2_nand2_2 U1679 (.A(keysched_new_key_o_84), .B(net24845), .Y(n1949));
sg13g2_inv_4 U1680 (.A(key_i_84_), .Y(n1948));
sg13g2_nand2_2 U1682 (.A(keysched_new_key_o_83), .B(net24837), .Y(n1951));
sg13g2_inv_4 U1683 (.A(key_i_83_), .Y(n1950));
sg13g2_nand2_2 U1685 (.A(keysched_new_key_o_82), .B(net24845), .Y(n1953));
sg13g2_inv_4 U1686 (.A(key_i_82_), .Y(n1952));
sg13g2_o21ai_1 U1687 (.A1(net26188), .A2(n1954), .B1(n1955), .Y(keysched_last_key_i_81));
sg13g2_nand2_2 U1688 (.A(keysched_new_key_o_81), .B(net25895), .Y(n1955));
sg13g2_inv_4 U1689 (.A(key_i_81_), .Y(n1954));
sg13g2_o21ai_1 U1690 (.A1(net26188), .A2(n1956), .B1(n1957), .Y(keysched_last_key_i_80));
sg13g2_nand2_2 U1691 (.A(keysched_new_key_o_80), .B(net25895), .Y(n1957));
sg13g2_inv_4 U1692 (.A(key_i_80_), .Y(n1956));
sg13g2_inv_4 U1695 (.A(key_i_7_), .Y(n862));
sg13g2_o21ai_1 U1696 (.A1(net24791), .A2(n1959), .B1(n1960), .Y(keysched_last_key_i_79));
sg13g2_nand2_2 U1697 (.A(keysched_new_key_o_79), .B(net25895), .Y(n1960));
sg13g2_inv_4 U1698 (.A(key_i_79_), .Y(n1959));
sg13g2_o21ai_1 U1699 (.A1(net26188), .A2(n1961), .B1(n1962), .Y(keysched_last_key_i_78));
sg13g2_nand2_2 U1700 (.A(keysched_new_key_o_78), .B(net25892), .Y(n1962));
sg13g2_inv_4 U1701 (.A(key_i_78_), .Y(n1961));
sg13g2_nand2_2 U1703 (.A(keysched_new_key_o_77), .B(net25892), .Y(n1964));
sg13g2_inv_4 U1704 (.A(key_i_77_), .Y(n1963));
sg13g2_o21ai_1 U1705 (.A1(net26188), .A2(n1965), .B1(n1966), .Y(keysched_last_key_i_76));
sg13g2_nand2_2 U1706 (.A(keysched_new_key_o_76), .B(net25895), .Y(n1966));
sg13g2_inv_4 U1707 (.A(key_i_76_), .Y(n1965));
sg13g2_nand2_2 U1709 (.A(keysched_new_key_o_75), .B(net24837), .Y(n1968));
sg13g2_inv_4 U1710 (.A(key_i_75_), .Y(n1967));
sg13g2_o21ai_1 U1711 (.A1(n4221), .A2(n1969), .B1(n1970), .Y(keysched_last_key_i_74));
sg13g2_nand2_2 U1712 (.A(keysched_new_key_o_74), .B(net24837), .Y(n1970));
sg13g2_inv_4 U1713 (.A(key_i_74_), .Y(n1969));
sg13g2_nand2_2 U1715 (.A(keysched_new_key_o_73), .B(net24837), .Y(n1972));
sg13g2_inv_4 U1716 (.A(key_i_73_), .Y(n1971));
sg13g2_o21ai_1 U1717 (.A1(net24801), .A2(n1973), .B1(n1974), .Y(keysched_last_key_i_72));
sg13g2_nand2_2 U1718 (.A(keysched_new_key_o_72), .B(net24837), .Y(n1974));
sg13g2_inv_4 U1719 (.A(key_i_72_), .Y(n1973));
sg13g2_o21ai_1 U1720 (.A1(net26188), .A2(n1975), .B1(n1976), .Y(keysched_last_key_i_71));
sg13g2_nand2_2 U1721 (.A(keysched_new_key_o_71), .B(net25895), .Y(n1976));
sg13g2_inv_4 U1722 (.A(key_i_71_), .Y(n1975));
sg13g2_o21ai_1 U1723 (.A1(net24795), .A2(n1977), .B1(n1978), .Y(keysched_last_key_i_70));
sg13g2_nand2_2 U1724 (.A(keysched_new_key_o_70), .B(net24837), .Y(n1978));
sg13g2_inv_4 U1725 (.A(key_i_70_), .Y(n1977));
sg13g2_inv_4 U1728 (.A(key_i_6_), .Y(n866));
sg13g2_o21ai_1 U1729 (.A1(net26188), .A2(n1980), .B1(n1981), .Y(keysched_last_key_i_69));
sg13g2_nand2_2 U1730 (.A(keysched_new_key_o_69), .B(net25895), .Y(n1981));
sg13g2_inv_4 U1731 (.A(key_i_69_), .Y(n1980));
sg13g2_o21ai_1 U1732 (.A1(net24795), .A2(n1982), .B1(n1983), .Y(keysched_last_key_i_68));
sg13g2_nand2_2 U1733 (.A(keysched_new_key_o_68), .B(net24837), .Y(n1983));
sg13g2_inv_4 U1734 (.A(key_i_68_), .Y(n1982));
sg13g2_o21ai_1 U1735 (.A1(net24795), .A2(n1984), .B1(n1985), .Y(keysched_last_key_i_67));
sg13g2_nand2_2 U1736 (.A(keysched_new_key_o_67), .B(net25895), .Y(n1985));
sg13g2_inv_4 U1737 (.A(key_i_67_), .Y(n1984));
sg13g2_o21ai_1 U1738 (.A1(net26188), .A2(n1986), .B1(n1987), .Y(keysched_last_key_i_66));
sg13g2_nand2_2 U1739 (.A(keysched_new_key_o_66), .B(net25895), .Y(n1987));
sg13g2_inv_4 U1740 (.A(key_i_66_), .Y(n1986));
sg13g2_o21ai_1 U1741 (.A1(net26188), .A2(n1988), .B1(n1989), .Y(keysched_last_key_i_65));
sg13g2_nand2_2 U1742 (.A(keysched_new_key_o_65), .B(n4155), .Y(n1989));
sg13g2_inv_4 U1743 (.A(key_i_65_), .Y(n1988));
sg13g2_nand2_2 U1745 (.A(keysched_new_key_o_64), .B(net24857), .Y(n1991));
sg13g2_inv_4 U1746 (.A(key_i_64_), .Y(n1990));
sg13g2_o21ai_1 U1747 (.A1(net26188), .A2(n870), .B1(n1992), .Y(keysched_last_key_i_63));
sg13g2_nand2_2 U1748 (.A(keysched_new_key_o_63), .B(net24845), .Y(n1992));
sg13g2_inv_4 U1749 (.A(key_i_63_), .Y(n870));
sg13g2_o21ai_1 U1750 (.A1(n4221), .A2(n874), .B1(n1993), .Y(keysched_last_key_i_62));
sg13g2_nand2_2 U1751 (.A(keysched_new_key_o_62), .B(net24857), .Y(n1993));
sg13g2_inv_4 U1752 (.A(key_i_62_), .Y(n874));
sg13g2_nand2_2 U1754 (.A(keysched_new_key_o_61), .B(n4155), .Y(n1994));
sg13g2_inv_4 U1755 (.A(key_i_61_), .Y(n878));
sg13g2_nand2_2 U1757 (.A(keysched_new_key_o_60), .B(n4155), .Y(n1995));
sg13g2_inv_4 U1758 (.A(key_i_60_), .Y(n882));
sg13g2_inv_4 U1761 (.A(key_i_5_), .Y(n886));
sg13g2_o21ai_1 U1762 (.A1(net24801), .A2(n890), .B1(n1997), .Y(keysched_last_key_i_59));
sg13g2_nand2_2 U1763 (.A(keysched_new_key_o_59), .B(net24857), .Y(n1997));
sg13g2_inv_4 U1764 (.A(key_i_59_), .Y(n890));
sg13g2_o21ai_1 U1765 (.A1(net24795), .A2(n894), .B1(n1998), .Y(keysched_last_key_i_58));
sg13g2_nand2_2 U1766 (.A(keysched_new_key_o_58), .B(net24837), .Y(n1998));
sg13g2_inv_4 U1767 (.A(key_i_58_), .Y(n894));
sg13g2_o21ai_1 U1768 (.A1(net26188), .A2(n898), .B1(n1999), .Y(keysched_last_key_i_57));
sg13g2_nand2_2 U1769 (.A(keysched_new_key_o_57), .B(net25895), .Y(n1999));
sg13g2_inv_4 U1770 (.A(key_i_57_), .Y(n898));
sg13g2_o21ai_1 U1771 (.A1(n4221), .A2(n902), .B1(n2000), .Y(keysched_last_key_i_56));
sg13g2_nand2_2 U1772 (.A(keysched_new_key_o_56), .B(n4156), .Y(n2000));
sg13g2_inv_4 U1773 (.A(key_i_56_), .Y(n902));
sg13g2_o21ai_1 U1774 (.A1(net24795), .A2(n906), .B1(n2001), .Y(keysched_last_key_i_55));
sg13g2_nand2_2 U1775 (.A(keysched_new_key_o_55), .B(net24837), .Y(n2001));
sg13g2_inv_4 U1776 (.A(key_i_55_), .Y(n906));
sg13g2_o21ai_1 U1777 (.A1(n4221), .A2(n910), .B1(n2002), .Y(keysched_last_key_i_54));
sg13g2_nand2_2 U1778 (.A(keysched_new_key_o_54), .B(net25892), .Y(n2002));
sg13g2_inv_4 U1779 (.A(key_i_54_), .Y(n910));
sg13g2_o21ai_1 U1780 (.A1(net26188), .A2(n914), .B1(n2003), .Y(keysched_last_key_i_53));
sg13g2_nand2_2 U1781 (.A(keysched_new_key_o_53), .B(net24837), .Y(n2003));
sg13g2_inv_4 U1782 (.A(key_i_53_), .Y(n914));
sg13g2_o21ai_1 U1783 (.A1(n4221), .A2(n918), .B1(n2004), .Y(keysched_last_key_i_52));
sg13g2_nand2_2 U1784 (.A(keysched_new_key_o_52), .B(net25895), .Y(n2004));
sg13g2_inv_4 U1785 (.A(key_i_52_), .Y(n918));
sg13g2_o21ai_1 U1786 (.A1(net26188), .A2(n922), .B1(n2005), .Y(keysched_last_key_i_51));
sg13g2_nand2_2 U1787 (.A(keysched_new_key_o_51), .B(net24837), .Y(n2005));
sg13g2_inv_4 U1788 (.A(key_i_51_), .Y(n922));
sg13g2_o21ai_1 U1789 (.A1(net26188), .A2(n926), .B1(n2006), .Y(keysched_last_key_i_50));
sg13g2_nand2_2 U1790 (.A(keysched_new_key_o_50), .B(net24837), .Y(n2006));
sg13g2_inv_4 U1791 (.A(key_i_50_), .Y(n926));
sg13g2_inv_4 U1794 (.A(key_i_4_), .Y(n930));
sg13g2_o21ai_1 U1795 (.A1(n4221), .A2(n934), .B1(n2008), .Y(keysched_last_key_i_49));
sg13g2_nand2_2 U1796 (.A(keysched_new_key_o_49), .B(net25895), .Y(n2008));
sg13g2_inv_4 U1797 (.A(key_i_49_), .Y(n934));
sg13g2_o21ai_1 U1798 (.A1(net24795), .A2(n938), .B1(n2009), .Y(keysched_last_key_i_48));
sg13g2_nand2_2 U1799 (.A(keysched_new_key_o_48), .B(net24837), .Y(n2009));
sg13g2_inv_4 U1800 (.A(key_i_48_), .Y(n938));
sg13g2_o21ai_1 U1801 (.A1(net26188), .A2(n942), .B1(n2010), .Y(keysched_last_key_i_47));
sg13g2_nand2_2 U1802 (.A(keysched_new_key_o_47), .B(net25895), .Y(n2010));
sg13g2_inv_4 U1803 (.A(key_i_47_), .Y(n942));
sg13g2_o21ai_1 U1804 (.A1(net26188), .A2(n946), .B1(n2011), .Y(keysched_last_key_i_46));
sg13g2_nand2_2 U1805 (.A(keysched_new_key_o_46), .B(net24837), .Y(n2011));
sg13g2_inv_4 U1806 (.A(key_i_46_), .Y(n946));
sg13g2_nand2_2 U1808 (.A(keysched_new_key_o_45), .B(net24837), .Y(n2012));
sg13g2_inv_4 U1809 (.A(key_i_45_), .Y(n950));
sg13g2_o21ai_1 U1810 (.A1(net24795), .A2(n954), .B1(n2013), .Y(keysched_last_key_i_44));
sg13g2_nand2_2 U1811 (.A(keysched_new_key_o_44), .B(net24837), .Y(n2013));
sg13g2_inv_4 U1812 (.A(key_i_44_), .Y(n954));
sg13g2_o21ai_1 U1813 (.A1(n4221), .A2(n958), .B1(n2014), .Y(keysched_last_key_i_43));
sg13g2_nand2_2 U1814 (.A(keysched_new_key_o_43), .B(net25895), .Y(n2014));
sg13g2_inv_4 U1815 (.A(key_i_43_), .Y(n958));
sg13g2_o21ai_1 U1816 (.A1(net24795), .A2(n962), .B1(n2015), .Y(keysched_last_key_i_42));
sg13g2_nand2_2 U1817 (.A(keysched_new_key_o_42), .B(net24837), .Y(n2015));
sg13g2_inv_4 U1818 (.A(key_i_42_), .Y(n962));
sg13g2_nand2_2 U1820 (.A(keysched_new_key_o_41), .B(net25895), .Y(n2016));
sg13g2_inv_4 U1821 (.A(key_i_41_), .Y(n966));
sg13g2_o21ai_1 U1822 (.A1(net26188), .A2(n970), .B1(n2017), .Y(keysched_last_key_i_40));
sg13g2_nand2_2 U1823 (.A(keysched_new_key_o_40), .B(net25895), .Y(n2017));
sg13g2_inv_4 U1824 (.A(key_i_40_), .Y(n970));
sg13g2_inv_4 U1827 (.A(key_i_3_), .Y(n974));
sg13g2_o21ai_1 U1828 (.A1(net24795), .A2(n978), .B1(n2019), .Y(keysched_last_key_i_39));
sg13g2_nand2_2 U1829 (.A(keysched_new_key_o_39), .B(net25895), .Y(n2019));
sg13g2_inv_4 U1830 (.A(key_i_39_), .Y(n978));
sg13g2_o21ai_1 U1831 (.A1(net26188), .A2(n982), .B1(n2020), .Y(keysched_last_key_i_38));
sg13g2_nand2_2 U1832 (.A(net25895), .B(keysched_new_key_o_38), .Y(n2020));
sg13g2_inv_4 U1833 (.A(key_i_38_), .Y(n982));
sg13g2_o21ai_1 U1834 (.A1(net24791), .A2(n986), .B1(n2021), .Y(keysched_last_key_i_37));
sg13g2_nand2_2 U1835 (.A(keysched_new_key_o_37), .B(net25895), .Y(n2021));
sg13g2_inv_4 U1836 (.A(key_i_37_), .Y(n986));
sg13g2_o21ai_1 U1837 (.A1(net24783), .A2(n990), .B1(n2022), .Y(keysched_last_key_i_36));
sg13g2_nand2_2 U1838 (.A(keysched_new_key_o_36), .B(net25895), .Y(n2022));
sg13g2_inv_4 U1839 (.A(key_i_36_), .Y(n990));
sg13g2_o21ai_1 U1840 (.A1(net24791), .A2(n994), .B1(n2023), .Y(keysched_last_key_i_35));
sg13g2_nand2_2 U1841 (.A(keysched_new_key_o_35), .B(n4155), .Y(n2023));
sg13g2_inv_4 U1842 (.A(key_i_35_), .Y(n994));
sg13g2_o21ai_1 U1843 (.A1(n4221), .A2(n998), .B1(n2024), .Y(keysched_last_key_i_34));
sg13g2_nand2_2 U1844 (.A(keysched_new_key_o_34), .B(net24847), .Y(n2024));
sg13g2_inv_4 U1845 (.A(key_i_34_), .Y(n998));
sg13g2_o21ai_1 U1846 (.A1(net24795), .A2(n1002), .B1(n2025), .Y(keysched_last_key_i_33));
sg13g2_nand2_2 U1847 (.A(keysched_new_key_o_33), .B(net25892), .Y(n2025));
sg13g2_inv_4 U1848 (.A(key_i_33_), .Y(n1002));
sg13g2_o21ai_1 U1849 (.A1(n4221), .A2(n1006), .B1(n2026), .Y(keysched_last_key_i_32));
sg13g2_nand2_2 U1850 (.A(keysched_new_key_o_32), .B(net25895), .Y(n2026));
sg13g2_inv_4 U1851 (.A(key_i_32_), .Y(n1006));
sg13g2_inv_4 U1854 (.A(key_i_31_), .Y(n1010));
sg13g2_inv_4 U1857 (.A(key_i_30_), .Y(n1014));
sg13g2_inv_4 U1860 (.A(key_i_2_), .Y(n1018));
sg13g2_inv_4 U1863 (.A(key_i_29_), .Y(n1022));
sg13g2_inv_4 U1866 (.A(key_i_28_), .Y(n1026));
sg13g2_inv_4 U1869 (.A(key_i_27_), .Y(n1030));
sg13g2_inv_4 U1872 (.A(key_i_26_), .Y(n1034));
sg13g2_inv_4 U1875 (.A(key_i_25_), .Y(n1038));
sg13g2_inv_4 U1878 (.A(key_i_24_), .Y(n1042));
sg13g2_inv_4 U1881 (.A(key_i_23_), .Y(n1046));
sg13g2_inv_4 U1884 (.A(key_i_22_), .Y(n1050));
sg13g2_inv_4 U1887 (.A(key_i_21_), .Y(n1054));
sg13g2_inv_4 U1890 (.A(key_i_20_), .Y(n1058));
sg13g2_inv_4 U1893 (.A(key_i_1_), .Y(n1062));
sg13g2_inv_4 U1896 (.A(key_i_19_), .Y(n1066));
sg13g2_inv_4 U1899 (.A(key_i_191_), .Y(n2042));
sg13g2_o21ai_1 U1900 (.A1(net24783), .A2(n2044), .B1(n2045), .Y(keysched_last_key_i_190));
sg13g2_nand2_2 U1901 (.A(keysched_new_key_o_190), .B(net24845), .Y(n2045));
sg13g2_inv_4 U1902 (.A(key_i_190_), .Y(n2044));
sg13g2_nand2_2 U1904 (.A(keysched_new_key_o_18), .B(net24847), .Y(n2046));
sg13g2_inv_4 U1905 (.A(key_i_18_), .Y(n1070));
sg13g2_nand2_2 U1907 (.A(keysched_new_key_o_189), .B(net24851), .Y(n2048));
sg13g2_inv_4 U1908 (.A(key_i_189_), .Y(n2047));
sg13g2_inv_4 U1911 (.A(key_i_188_), .Y(n2049));
sg13g2_nand2_2 U1913 (.A(keysched_new_key_o_187), .B(net25895), .Y(n2052));
sg13g2_inv_4 U1914 (.A(key_i_187_), .Y(n2051));
sg13g2_nand2_2 U1916 (.A(keysched_new_key_o_186), .B(net24857), .Y(n2054));
sg13g2_inv_4 U1917 (.A(key_i_186_), .Y(n2053));
sg13g2_nand2_2 U1919 (.A(keysched_new_key_o_185), .B(net25895), .Y(n2056));
sg13g2_inv_4 U1920 (.A(key_i_185_), .Y(n2055));
sg13g2_nand2_2 U1922 (.A(keysched_new_key_o_184), .B(n4156), .Y(n2058));
sg13g2_inv_4 U1923 (.A(key_i_184_), .Y(n2057));
sg13g2_inv_4 U1926 (.A(key_i_183_), .Y(n2059));
sg13g2_o21ai_1 U1927 (.A1(net24791), .A2(n2061), .B1(n2062), .Y(keysched_last_key_i_182));
sg13g2_nand2_2 U1928 (.A(keysched_new_key_o_182), .B(net24845), .Y(n2062));
sg13g2_inv_4 U1929 (.A(key_i_182_), .Y(n2061));
sg13g2_nand2_2 U1931 (.A(keysched_new_key_o_181), .B(net24851), .Y(n2064));
sg13g2_inv_4 U1932 (.A(key_i_181_), .Y(n2063));
sg13g2_nand2_2 U1934 (.A(keysched_new_key_o_180), .B(net24857), .Y(n2066));
sg13g2_inv_4 U1935 (.A(key_i_180_), .Y(n2065));
sg13g2_inv_4 U1938 (.A(key_i_17_), .Y(n1074));
sg13g2_nand2_2 U1940 (.A(keysched_new_key_o_179), .B(net24837), .Y(n2069));
sg13g2_inv_4 U1941 (.A(key_i_179_), .Y(n2068));
sg13g2_o21ai_1 U1942 (.A1(net24791), .A2(n2070), .B1(n2071), .Y(keysched_last_key_i_178));
sg13g2_nand2_2 U1943 (.A(keysched_new_key_o_178), .B(net24837), .Y(n2071));
sg13g2_inv_4 U1944 (.A(key_i_178_), .Y(n2070));
sg13g2_nand2_2 U1946 (.A(keysched_new_key_o_177), .B(net24837), .Y(n2073));
sg13g2_inv_4 U1947 (.A(key_i_177_), .Y(n2072));
sg13g2_nand2_2 U1949 (.A(keysched_new_key_o_176), .B(net24837), .Y(n2075));
sg13g2_inv_4 U1950 (.A(key_i_176_), .Y(n2074));
sg13g2_nand2_2 U1952 (.A(keysched_new_key_o_175), .B(net24837), .Y(n2077));
sg13g2_inv_4 U1953 (.A(key_i_175_), .Y(n2076));
sg13g2_o21ai_1 U1954 (.A1(net24791), .A2(n2078), .B1(n2079), .Y(keysched_last_key_i_174));
sg13g2_nand2_2 U1955 (.A(keysched_new_key_o_174), .B(net25892), .Y(n2079));
sg13g2_inv_4 U1956 (.A(key_i_174_), .Y(n2078));
sg13g2_o21ai_1 U1957 (.A1(net24791), .A2(n2080), .B1(n2081), .Y(keysched_last_key_i_173));
sg13g2_nand2_2 U1958 (.A(keysched_new_key_o_173), .B(net25892), .Y(n2081));
sg13g2_inv_4 U1959 (.A(key_i_173_), .Y(n2080));
sg13g2_nand2_2 U1961 (.A(keysched_new_key_o_172), .B(net24845), .Y(n2083));
sg13g2_inv_4 U1962 (.A(key_i_172_), .Y(n2082));
sg13g2_o21ai_1 U1963 (.A1(net24791), .A2(n2084), .B1(n2085), .Y(keysched_last_key_i_171));
sg13g2_nand2_2 U1964 (.A(keysched_new_key_o_171), .B(net25892), .Y(n2085));
sg13g2_inv_4 U1965 (.A(key_i_171_), .Y(n2084));
sg13g2_o21ai_1 U1966 (.A1(net24791), .A2(n2086), .B1(n2087), .Y(keysched_last_key_i_170));
sg13g2_nand2_2 U1967 (.A(keysched_new_key_o_170), .B(net25892), .Y(n2087));
sg13g2_inv_4 U1968 (.A(key_i_170_), .Y(n2086));
sg13g2_inv_4 U1971 (.A(key_i_16_), .Y(n1078));
sg13g2_o21ai_1 U1972 (.A1(net26188), .A2(n2089), .B1(n2090), .Y(keysched_last_key_i_169));
sg13g2_nand2_2 U1973 (.A(keysched_new_key_o_169), .B(net24845), .Y(n2090));
sg13g2_inv_4 U1974 (.A(key_i_169_), .Y(n2089));
sg13g2_nand2_2 U1976 (.A(keysched_new_key_o_168), .B(net25895), .Y(n2092));
sg13g2_inv_4 U1977 (.A(key_i_168_), .Y(n2091));
sg13g2_nand2_2 U1979 (.A(keysched_new_key_o_167), .B(net25895), .Y(n2094));
sg13g2_inv_4 U1980 (.A(key_i_167_), .Y(n2093));
sg13g2_nand2_2 U1982 (.A(keysched_new_key_o_166), .B(net25895), .Y(n2096));
sg13g2_inv_4 U1983 (.A(key_i_166_), .Y(n2095));
sg13g2_nand2_2 U1985 (.A(keysched_new_key_o_165), .B(net25895), .Y(n2098));
sg13g2_inv_4 U1986 (.A(key_i_165_), .Y(n2097));
sg13g2_nand2_2 U1988 (.A(keysched_new_key_o_164), .B(net25895), .Y(n2100));
sg13g2_inv_4 U1989 (.A(key_i_164_), .Y(n2099));
sg13g2_o21ai_1 U1990 (.A1(net24795), .A2(n2101), .B1(n2102), .Y(keysched_last_key_i_163));
sg13g2_nand2_2 U1991 (.A(keysched_new_key_o_163), .B(net25895), .Y(n2102));
sg13g2_inv_4 U1992 (.A(key_i_163_), .Y(n2101));
sg13g2_o21ai_1 U1993 (.A1(net24795), .A2(n2103), .B1(n2104), .Y(keysched_last_key_i_162));
sg13g2_nand2_2 U1994 (.A(keysched_new_key_o_162), .B(net25895), .Y(n2104));
sg13g2_inv_4 U1995 (.A(key_i_162_), .Y(n2103));
sg13g2_nand2_2 U1997 (.A(keysched_new_key_o_161), .B(net25895), .Y(n2106));
sg13g2_inv_4 U1998 (.A(key_i_161_), .Y(n2105));
sg13g2_nand2_2 U2000 (.A(keysched_new_key_o_160), .B(net25895), .Y(n2108));
sg13g2_inv_4 U2001 (.A(key_i_160_), .Y(n2107));
sg13g2_nand2_2 U2006 (.A(keysched_new_key_o_159), .B(net24837), .Y(n2111));
sg13g2_inv_4 U2007 (.A(key_i_159_), .Y(n2110));
sg13g2_o21ai_1 U2008 (.A1(net24783), .A2(n2112), .B1(n2113), .Y(keysched_last_key_i_158));
sg13g2_nand2_2 U2009 (.A(keysched_new_key_o_158), .B(net24837), .Y(n2113));
sg13g2_inv_4 U2010 (.A(key_i_158_), .Y(n2112));
sg13g2_o21ai_1 U2011 (.A1(net24801), .A2(n2114), .B1(n2115), .Y(keysched_last_key_i_157));
sg13g2_nand2_2 U2012 (.A(keysched_new_key_o_157), .B(net24837), .Y(n2115));
sg13g2_inv_4 U2013 (.A(key_i_157_), .Y(n2114));
sg13g2_o21ai_1 U2014 (.A1(net24801), .A2(n2116), .B1(n2117), .Y(keysched_last_key_i_156));
sg13g2_nand2_2 U2015 (.A(keysched_new_key_o_156), .B(net24837), .Y(n2117));
sg13g2_inv_4 U2016 (.A(key_i_156_), .Y(n2116));
sg13g2_o21ai_1 U2017 (.A1(net24783), .A2(n2118), .B1(n2119), .Y(keysched_last_key_i_155));
sg13g2_nand2_2 U2018 (.A(keysched_new_key_o_155), .B(net24837), .Y(n2119));
sg13g2_inv_4 U2019 (.A(key_i_155_), .Y(n2118));
sg13g2_o21ai_1 U2020 (.A1(net26188), .A2(n2120), .B1(n2121), .Y(keysched_last_key_i_154));
sg13g2_nand2_2 U2021 (.A(keysched_new_key_o_154), .B(net24837), .Y(n2121));
sg13g2_inv_4 U2022 (.A(key_i_154_), .Y(n2120));
sg13g2_o21ai_1 U2023 (.A1(net24783), .A2(n2122), .B1(n2123), .Y(keysched_last_key_i_153));
sg13g2_nand2_2 U2024 (.A(keysched_new_key_o_153), .B(net24837), .Y(n2123));
sg13g2_inv_4 U2025 (.A(key_i_153_), .Y(n2122));
sg13g2_o21ai_1 U2026 (.A1(net24801), .A2(n2124), .B1(n2125), .Y(keysched_last_key_i_152));
sg13g2_nand2_2 U2027 (.A(keysched_new_key_o_152), .B(net24837), .Y(n2125));
sg13g2_inv_4 U2028 (.A(key_i_152_), .Y(n2124));
sg13g2_o21ai_1 U2029 (.A1(net24795), .A2(n2126), .B1(n2127), .Y(keysched_last_key_i_151));
sg13g2_nand2_2 U2030 (.A(keysched_new_key_o_151), .B(net24837), .Y(n2127));
sg13g2_inv_4 U2031 (.A(key_i_151_), .Y(n2126));
sg13g2_o21ai_1 U2032 (.A1(net24783), .A2(n2128), .B1(n2129), .Y(keysched_last_key_i_150));
sg13g2_nand2_2 U2033 (.A(keysched_new_key_o_150), .B(net24837), .Y(n2129));
sg13g2_inv_4 U2034 (.A(key_i_150_), .Y(n2128));
sg13g2_inv_4 U2037 (.A(key_i_14_), .Y(n1086));
sg13g2_o21ai_1 U2038 (.A1(net24791), .A2(n2131), .B1(n2132), .Y(keysched_last_key_i_149));
sg13g2_nand2_2 U2039 (.A(keysched_new_key_o_149), .B(net24837), .Y(n2132));
sg13g2_inv_4 U2040 (.A(key_i_149_), .Y(n2131));
sg13g2_o21ai_1 U2041 (.A1(n4221), .A2(n2133), .B1(n2134), .Y(keysched_last_key_i_148));
sg13g2_nand2_2 U2042 (.A(keysched_new_key_o_148), .B(net25895), .Y(n2134));
sg13g2_inv_4 U2043 (.A(key_i_148_), .Y(n2133));
sg13g2_nand2_2 U2045 (.A(keysched_new_key_o_147), .B(net25895), .Y(n2136));
sg13g2_inv_4 U2046 (.A(key_i_147_), .Y(n2135));
sg13g2_nand2_2 U2048 (.A(keysched_new_key_o_146), .B(net25895), .Y(n2138));
sg13g2_inv_4 U2049 (.A(key_i_146_), .Y(n2137));
sg13g2_nand2_2 U2051 (.A(keysched_new_key_o_145), .B(net25895), .Y(n2140));
sg13g2_inv_4 U2052 (.A(key_i_145_), .Y(n2139));
sg13g2_o21ai_1 U2053 (.A1(net26188), .A2(n2141), .B1(n2142), .Y(keysched_last_key_i_144));
sg13g2_nand2_2 U2054 (.A(keysched_new_key_o_144), .B(net25895), .Y(n2142));
sg13g2_inv_4 U2055 (.A(key_i_144_), .Y(n2141));
sg13g2_o21ai_1 U2056 (.A1(net26188), .A2(n2143), .B1(n2144), .Y(keysched_last_key_i_143));
sg13g2_nand2_2 U2057 (.A(keysched_new_key_o_143), .B(net25895), .Y(n2144));
sg13g2_inv_4 U2058 (.A(key_i_143_), .Y(n2143));
sg13g2_o21ai_1 U2059 (.A1(net24791), .A2(n2145), .B1(n2146), .Y(keysched_last_key_i_142));
sg13g2_nand2_2 U2060 (.A(keysched_new_key_o_142), .B(net24839), .Y(n2146));
sg13g2_inv_4 U2061 (.A(key_i_142_), .Y(n2145));
sg13g2_nand2_2 U2063 (.A(keysched_new_key_o_141), .B(net24839), .Y(n2148));
sg13g2_inv_4 U2064 (.A(key_i_141_), .Y(n2147));
sg13g2_o21ai_1 U2065 (.A1(net24795), .A2(n2149), .B1(n2150), .Y(keysched_last_key_i_140));
sg13g2_nand2_2 U2066 (.A(keysched_new_key_o_140), .B(net24837), .Y(n2150));
sg13g2_inv_4 U2067 (.A(key_i_140_), .Y(n2149));
sg13g2_inv_4 U2070 (.A(key_i_13_), .Y(n1090));
sg13g2_o21ai_1 U2071 (.A1(net24791), .A2(n2152), .B1(n2153), .Y(keysched_last_key_i_139));
sg13g2_nand2_2 U2072 (.A(keysched_new_key_o_139), .B(net24845), .Y(n2153));
sg13g2_inv_4 U2073 (.A(key_i_139_), .Y(n2152));
sg13g2_o21ai_1 U2074 (.A1(n4221), .A2(n2154), .B1(n2155), .Y(keysched_last_key_i_138));
sg13g2_nand2_2 U2075 (.A(keysched_new_key_o_138), .B(net24845), .Y(n2155));
sg13g2_inv_4 U2076 (.A(key_i_138_), .Y(n2154));
sg13g2_o21ai_1 U2077 (.A1(n4221), .A2(n2156), .B1(n2157), .Y(keysched_last_key_i_137));
sg13g2_nand2_2 U2078 (.A(keysched_new_key_o_137), .B(net24845), .Y(n2157));
sg13g2_inv_4 U2079 (.A(key_i_137_), .Y(n2156));
sg13g2_nand2_2 U2081 (.A(keysched_new_key_o_136), .B(net24837), .Y(n2159));
sg13g2_inv_4 U2082 (.A(key_i_136_), .Y(n2158));
sg13g2_o21ai_1 U2083 (.A1(net24795), .A2(n2160), .B1(n2161), .Y(keysched_last_key_i_135));
sg13g2_nand2_2 U2084 (.A(keysched_new_key_o_135), .B(net24845), .Y(n2161));
sg13g2_inv_4 U2085 (.A(key_i_135_), .Y(n2160));
sg13g2_o21ai_1 U2086 (.A1(net26188), .A2(n2162), .B1(n2163), .Y(keysched_last_key_i_134));
sg13g2_nand2_2 U2087 (.A(keysched_new_key_o_134), .B(net24837), .Y(n2163));
sg13g2_inv_4 U2088 (.A(key_i_134_), .Y(n2162));
sg13g2_o21ai_1 U2089 (.A1(n4221), .A2(n2164), .B1(n2165), .Y(keysched_last_key_i_133));
sg13g2_nand2_2 U2090 (.A(keysched_new_key_o_133), .B(net24837), .Y(n2165));
sg13g2_inv_4 U2091 (.A(key_i_133_), .Y(n2164));
sg13g2_o21ai_1 U2092 (.A1(net26188), .A2(n2166), .B1(n2167), .Y(keysched_last_key_i_132));
sg13g2_nand2_2 U2093 (.A(keysched_new_key_o_132), .B(net24845), .Y(n2167));
sg13g2_inv_4 U2094 (.A(key_i_132_), .Y(n2166));
sg13g2_o21ai_1 U2095 (.A1(n4221), .A2(n2168), .B1(n2169), .Y(keysched_last_key_i_131));
sg13g2_nand2_2 U2096 (.A(keysched_new_key_o_131), .B(net24845), .Y(n2169));
sg13g2_inv_4 U2097 (.A(key_i_131_), .Y(n2168));
sg13g2_o21ai_1 U2098 (.A1(net24795), .A2(n2170), .B1(n2171), .Y(keysched_last_key_i_130));
sg13g2_nand2_2 U2099 (.A(keysched_new_key_o_130), .B(net24837), .Y(n2171));
sg13g2_inv_4 U2100 (.A(key_i_130_), .Y(n2170));
sg13g2_inv_4 U2103 (.A(key_i_12_), .Y(n1094));
sg13g2_nand2_2 U2105 (.A(keysched_new_key_o_129), .B(net24837), .Y(n2174));
sg13g2_nand2_2 U2108 (.A(keysched_new_key_o_128), .B(net24837), .Y(n2176));
sg13g2_inv_4 U2109 (.A(key_i_128_), .Y(n2175));
sg13g2_o21ai_1 U2110 (.A1(net26188), .A2(n2177), .B1(n2178), .Y(keysched_last_key_i_127));
sg13g2_nand2_2 U2111 (.A(keysched_new_key_o_127), .B(net25892), .Y(n2178));
sg13g2_inv_4 U2112 (.A(key_i_127_), .Y(n2177));
sg13g2_o21ai_1 U2113 (.A1(net24795), .A2(n2179), .B1(n2180), .Y(keysched_last_key_i_126));
sg13g2_nand2_2 U2114 (.A(keysched_new_key_o_126), .B(net24837), .Y(n2180));
sg13g2_inv_4 U2115 (.A(key_i_126_), .Y(n2179));
sg13g2_o21ai_1 U2116 (.A1(net24783), .A2(n2181), .B1(n2182), .Y(keysched_last_key_i_125));
sg13g2_nand2_2 U2117 (.A(keysched_new_key_o_125), .B(net24845), .Y(n2182));
sg13g2_inv_4 U2118 (.A(key_i_125_), .Y(n2181));
sg13g2_o21ai_1 U2119 (.A1(net26188), .A2(n2183), .B1(n2184), .Y(keysched_last_key_i_124));
sg13g2_nand2_2 U2120 (.A(keysched_new_key_o_124), .B(net24845), .Y(n2184));
sg13g2_inv_4 U2121 (.A(key_i_124_), .Y(n2183));
sg13g2_o21ai_1 U2122 (.A1(net24801), .A2(n2185), .B1(n2186), .Y(keysched_last_key_i_123));
sg13g2_nand2_2 U2123 (.A(keysched_new_key_o_123), .B(net24837), .Y(n2186));
sg13g2_inv_4 U2124 (.A(key_i_123_), .Y(n2185));
sg13g2_o21ai_1 U2125 (.A1(net26188), .A2(n2187), .B1(n2188), .Y(keysched_last_key_i_122));
sg13g2_nand2_2 U2126 (.A(keysched_new_key_o_122), .B(net24837), .Y(n2188));
sg13g2_inv_4 U2127 (.A(key_i_122_), .Y(n2187));
sg13g2_o21ai_1 U2128 (.A1(net26188), .A2(n2189), .B1(n2190), .Y(keysched_last_key_i_121));
sg13g2_nand2_2 U2129 (.A(keysched_new_key_o_121), .B(net25892), .Y(n2190));
sg13g2_inv_4 U2130 (.A(key_i_121_), .Y(n2189));
sg13g2_o21ai_1 U2131 (.A1(net24783), .A2(n2191), .B1(n2192), .Y(keysched_last_key_i_120));
sg13g2_nand2_2 U2132 (.A(keysched_new_key_o_120), .B(net24837), .Y(n2192));
sg13g2_inv_4 U2133 (.A(key_i_120_), .Y(n2191));
sg13g2_inv_4 U2136 (.A(key_i_11_), .Y(n1098));
sg13g2_o21ai_1 U2137 (.A1(n4221), .A2(n2194), .B1(n2195), .Y(keysched_last_key_i_119));
sg13g2_nand2_2 U2138 (.A(keysched_new_key_o_119), .B(net25895), .Y(n2195));
sg13g2_inv_4 U2139 (.A(key_i_119_), .Y(n2194));
sg13g2_o21ai_1 U2140 (.A1(net26188), .A2(n2196), .B1(n2197), .Y(keysched_last_key_i_118));
sg13g2_nand2_2 U2141 (.A(keysched_new_key_o_118), .B(net25895), .Y(n2197));
sg13g2_inv_4 U2142 (.A(key_i_118_), .Y(n2196));
sg13g2_o21ai_1 U2143 (.A1(n4221), .A2(n2198), .B1(n2199), .Y(keysched_last_key_i_117));
sg13g2_nand2_2 U2144 (.A(keysched_new_key_o_117), .B(net25895), .Y(n2199));
sg13g2_inv_4 U2145 (.A(key_i_117_), .Y(n2198));
sg13g2_o21ai_1 U2146 (.A1(n4221), .A2(n2200), .B1(n2201), .Y(keysched_last_key_i_116));
sg13g2_nand2_2 U2147 (.A(keysched_new_key_o_116), .B(net25895), .Y(n2201));
sg13g2_inv_4 U2148 (.A(key_i_116_), .Y(n2200));
sg13g2_o21ai_1 U2149 (.A1(n4221), .A2(n2202), .B1(n2203), .Y(keysched_last_key_i_115));
sg13g2_nand2_2 U2150 (.A(keysched_new_key_o_115), .B(net25895), .Y(n2203));
sg13g2_inv_4 U2151 (.A(key_i_115_), .Y(n2202));
sg13g2_o21ai_1 U2152 (.A1(net24801), .A2(n2204), .B1(n2205), .Y(keysched_last_key_i_114));
sg13g2_nand2_2 U2153 (.A(keysched_new_key_o_114), .B(net25895), .Y(n2205));
sg13g2_inv_4 U2154 (.A(key_i_114_), .Y(n2204));
sg13g2_o21ai_1 U2155 (.A1(net26188), .A2(n2206), .B1(n2207), .Y(keysched_last_key_i_113));
sg13g2_nand2_2 U2156 (.A(keysched_new_key_o_113), .B(net25895), .Y(n2207));
sg13g2_inv_4 U2157 (.A(key_i_113_), .Y(n2206));
sg13g2_o21ai_1 U2158 (.A1(n4221), .A2(n2208), .B1(n2209), .Y(keysched_last_key_i_112));
sg13g2_nand2_2 U2159 (.A(keysched_new_key_o_112), .B(net25895), .Y(n2209));
sg13g2_inv_4 U2160 (.A(key_i_112_), .Y(n2208));
sg13g2_o21ai_1 U2161 (.A1(net26188), .A2(n2210), .B1(n2211), .Y(keysched_last_key_i_111));
sg13g2_nand2_2 U2162 (.A(keysched_new_key_o_111), .B(net25895), .Y(n2211));
sg13g2_inv_4 U2163 (.A(key_i_111_), .Y(n2210));
sg13g2_o21ai_1 U2164 (.A1(net26188), .A2(n2212), .B1(n2213), .Y(keysched_last_key_i_110));
sg13g2_nand2_2 U2165 (.A(keysched_new_key_o_110), .B(net24839), .Y(n2213));
sg13g2_inv_4 U2166 (.A(key_i_110_), .Y(n2212));
sg13g2_inv_4 U2169 (.A(key_i_10_), .Y(n1102));
sg13g2_o21ai_1 U2170 (.A1(net26188), .A2(n2215), .B1(n2216), .Y(keysched_last_key_i_109));
sg13g2_nand2_2 U2171 (.A(keysched_new_key_o_109), .B(net25895), .Y(n2216));
sg13g2_inv_4 U2172 (.A(key_i_109_), .Y(n2215));
sg13g2_o21ai_1 U2173 (.A1(net24795), .A2(n2217), .B1(n2218), .Y(keysched_last_key_i_108));
sg13g2_nand2_2 U2174 (.A(keysched_new_key_o_108), .B(net25895), .Y(n2218));
sg13g2_inv_4 U2175 (.A(key_i_108_), .Y(n2217));
sg13g2_o21ai_1 U2176 (.A1(net24791), .A2(n2219), .B1(n2220), .Y(keysched_last_key_i_107));
sg13g2_nand2_2 U2177 (.A(keysched_new_key_o_107), .B(net25895), .Y(n2220));
sg13g2_inv_4 U2178 (.A(key_i_107_), .Y(n2219));
sg13g2_nand2_2 U2180 (.A(keysched_new_key_o_106), .B(net25895), .Y(n2222));
sg13g2_inv_4 U2181 (.A(key_i_106_), .Y(n2221));
sg13g2_nand2_2 U2183 (.A(keysched_new_key_o_105), .B(net25895), .Y(n2224));
sg13g2_inv_4 U2184 (.A(key_i_105_), .Y(n2223));
sg13g2_nand2_2 U2186 (.A(keysched_new_key_o_104), .B(net25895), .Y(n2226));
sg13g2_inv_4 U2187 (.A(key_i_104_), .Y(n2225));
sg13g2_o21ai_1 U2188 (.A1(net26188), .A2(n2227), .B1(n2228), .Y(keysched_last_key_i_103));
sg13g2_nand2_2 U2189 (.A(keysched_new_key_o_103), .B(net25895), .Y(n2228));
sg13g2_inv_4 U2190 (.A(key_i_103_), .Y(n2227));
sg13g2_nand2_2 U2192 (.A(keysched_new_key_o_102), .B(net25895), .Y(n2230));
sg13g2_inv_4 U2193 (.A(key_i_102_), .Y(n2229));
sg13g2_nand2_2 U2195 (.A(keysched_new_key_o_101), .B(net25895), .Y(n2232));
sg13g2_inv_4 U2196 (.A(key_i_101_), .Y(n2231));
sg13g2_nand2_2 U2198 (.A(keysched_new_key_o_100), .B(net25895), .Y(n2234));
sg13g2_inv_4 U2199 (.A(key_i_100_), .Y(n2233));
sg13g2_inv_4 U2205 (.A(keysched_ready_o), .Y(n1131));
sg13g2_inv_4 U2206 (.A(key_i_0_), .Y(n1106));
sg13g2_a21oi_2 U2224 (.A1(n2244), .A2(n2245), .B1(n2246), .Y(n2243));
sg13g2_nor2_2 U2225 (.A(n2247), .B(n2248), .Y(n2246));
sg13g2_o21ai_1 U2226 (.A1(n4167), .A2(n2247), .B1(n2249), .Y(n2245));
sg13g2_a21oi_2 U2227 (.A1(n4315), .A2(n2250), .B1(n2251), .Y(n2249));
sg13g2_nor2_2 U2228 (.A(n4165), .B(n558), .Y(n2251));
sg13g2_inv_4 U2229 (.A(n2250), .Y(n2242));
sg13g2_o21ai_1 U2230 (.A1(n4329), .A2(n2247), .B1(n2252), .Y(n2250));
sg13g2_a21oi_2 U2231 (.A1(data_i_9_), .A2(n4307), .B1(n2254), .Y(n2252));
sg13g2_nor2_2 U2232 (.A(n555), .B(n558), .Y(n2254));
sg13g2_inv_4 U2233 (.A(mixcol_data_o_9), .Y(n558));
sg13g2_inv_4 U2234 (.A(subbytes_data_o_9), .Y(n2247));
sg13g2_a21oi_2 U2236 (.A1(n2244), .A2(n2257), .B1(n2258), .Y(n2256));
sg13g2_nor2_2 U2237 (.A(n2259), .B(n2248), .Y(n2258));
sg13g2_o21ai_1 U2238 (.A1(n553), .A2(n2259), .B1(n2260), .Y(n2257));
sg13g2_a21oi_2 U2239 (.A1(n4315), .A2(n2261), .B1(n2262), .Y(n2260));
sg13g2_nor2_2 U2240 (.A(n4164), .B(n561), .Y(n2262));
sg13g2_inv_4 U2241 (.A(n2261), .Y(n2255));
sg13g2_o21ai_1 U2242 (.A1(n4327), .A2(n2259), .B1(n2263), .Y(n2261));
sg13g2_a21oi_2 U2243 (.A1(data_i_99_), .A2(n4307), .B1(n2264), .Y(n2263));
sg13g2_nor2_2 U2244 (.A(n555), .B(n561), .Y(n2264));
sg13g2_inv_4 U2245 (.A(mixcol_data_o_99), .Y(n561));
sg13g2_inv_4 U2246 (.A(subbytes_data_o_99), .Y(n2259));
sg13g2_a21oi_2 U2248 (.A1(n4313), .A2(n2267), .B1(n2268), .Y(n2266));
sg13g2_nor2_2 U2249 (.A(n2269), .B(n2248), .Y(n2268));
sg13g2_o21ai_1 U2250 (.A1(n4167), .A2(n2269), .B1(n2270), .Y(n2267));
sg13g2_a21oi_2 U2251 (.A1(n4315), .A2(n2271), .B1(n2272), .Y(n2270));
sg13g2_nor2_2 U2252 (.A(n4165), .B(n563), .Y(n2272));
sg13g2_inv_4 U2253 (.A(n2271), .Y(n2265));
sg13g2_o21ai_1 U2254 (.A1(n4326), .A2(n2269), .B1(n2273), .Y(n2271));
sg13g2_a21oi_2 U2255 (.A1(data_i_98_), .A2(n4308), .B1(n2274), .Y(n2273));
sg13g2_nor2_2 U2256 (.A(n555), .B(n563), .Y(n2274));
sg13g2_inv_4 U2257 (.A(mixcol_data_o_98), .Y(n563));
sg13g2_inv_4 U2258 (.A(subbytes_data_o_98), .Y(n2269));
sg13g2_a21oi_2 U2260 (.A1(n4312), .A2(n2277), .B1(n2278), .Y(n2276));
sg13g2_nor2_2 U2261 (.A(n2279), .B(n2248), .Y(n2278));
sg13g2_o21ai_1 U2262 (.A1(n553), .A2(n2279), .B1(n2280), .Y(n2277));
sg13g2_a21oi_2 U2263 (.A1(n4315), .A2(n2281), .B1(n2282), .Y(n2280));
sg13g2_nor2_2 U2264 (.A(n4165), .B(n565), .Y(n2282));
sg13g2_inv_4 U2265 (.A(n2281), .Y(n2275));
sg13g2_o21ai_1 U2266 (.A1(n4325), .A2(n2279), .B1(n2283), .Y(n2281));
sg13g2_a21oi_2 U2267 (.A1(data_i_97_), .A2(n4308), .B1(n2284), .Y(n2283));
sg13g2_nor2_2 U2268 (.A(n555), .B(n565), .Y(n2284));
sg13g2_inv_4 U2269 (.A(mixcol_data_o_97), .Y(n565));
sg13g2_inv_4 U2270 (.A(subbytes_data_o_97), .Y(n2279));
sg13g2_a21oi_2 U2272 (.A1(n2244), .A2(n2287), .B1(n2288), .Y(n2286));
sg13g2_nor2_2 U2273 (.A(n2289), .B(n2248), .Y(n2288));
sg13g2_o21ai_1 U2274 (.A1(n4167), .A2(n2289), .B1(n2290), .Y(n2287));
sg13g2_a21oi_2 U2275 (.A1(n4315), .A2(n2291), .B1(n2292), .Y(n2290));
sg13g2_nor2_2 U2276 (.A(n4164), .B(n567), .Y(n2292));
sg13g2_inv_4 U2277 (.A(n2291), .Y(n2285));
sg13g2_o21ai_1 U2278 (.A1(n4330), .A2(n2289), .B1(n2293), .Y(n2291));
sg13g2_a21oi_2 U2279 (.A1(data_i_96_), .A2(n4308), .B1(n2294), .Y(n2293));
sg13g2_nor2_2 U2280 (.A(n555), .B(n567), .Y(n2294));
sg13g2_inv_4 U2281 (.A(mixcol_data_o_96), .Y(n567));
sg13g2_inv_4 U2282 (.A(subbytes_data_o_96), .Y(n2289));
sg13g2_a21oi_2 U2284 (.A1(n4313), .A2(n2297), .B1(n2298), .Y(n2296));
sg13g2_nor2_2 U2285 (.A(n2299), .B(n2248), .Y(n2298));
sg13g2_o21ai_1 U2286 (.A1(n553), .A2(n2299), .B1(n2300), .Y(n2297));
sg13g2_a21oi_2 U2287 (.A1(n4315), .A2(n2301), .B1(n2302), .Y(n2300));
sg13g2_nor2_2 U2288 (.A(n4165), .B(n569), .Y(n2302));
sg13g2_inv_4 U2289 (.A(n2301), .Y(n2295));
sg13g2_o21ai_1 U2290 (.A1(n4328), .A2(n2299), .B1(n2303), .Y(n2301));
sg13g2_a21oi_2 U2291 (.A1(data_i_95_), .A2(n4308), .B1(n2304), .Y(n2303));
sg13g2_nor2_2 U2292 (.A(n555), .B(n569), .Y(n2304));
sg13g2_inv_4 U2293 (.A(mixcol_data_o_95), .Y(n569));
sg13g2_inv_4 U2294 (.A(subbytes_data_o_95), .Y(n2299));
sg13g2_a21oi_2 U2296 (.A1(n4312), .A2(n2307), .B1(n2308), .Y(n2306));
sg13g2_nor2_2 U2297 (.A(n2309), .B(n2248), .Y(n2308));
sg13g2_o21ai_1 U2298 (.A1(n4167), .A2(n2309), .B1(n2310), .Y(n2307));
sg13g2_a21oi_2 U2299 (.A1(n4315), .A2(n2311), .B1(n2312), .Y(n2310));
sg13g2_nor2_2 U2300 (.A(n4164), .B(n571), .Y(n2312));
sg13g2_inv_4 U2301 (.A(n2311), .Y(n2305));
sg13g2_o21ai_1 U2302 (.A1(n4329), .A2(n2309), .B1(n2313), .Y(n2311));
sg13g2_a21oi_2 U2303 (.A1(data_i_94_), .A2(n4308), .B1(n2314), .Y(n2313));
sg13g2_nor2_2 U2304 (.A(n555), .B(n571), .Y(n2314));
sg13g2_inv_4 U2305 (.A(mixcol_data_o_94), .Y(n571));
sg13g2_inv_4 U2306 (.A(subbytes_data_o_94), .Y(n2309));
sg13g2_a21oi_2 U2308 (.A1(n4312), .A2(n2317), .B1(n2318), .Y(n2316));
sg13g2_nor2_2 U2309 (.A(n2319), .B(n2248), .Y(n2318));
sg13g2_o21ai_1 U2310 (.A1(n4167), .A2(n2319), .B1(n2320), .Y(n2317));
sg13g2_a21oi_2 U2311 (.A1(n4315), .A2(n2321), .B1(n2322), .Y(n2320));
sg13g2_nor2_2 U2312 (.A(n4164), .B(n573), .Y(n2322));
sg13g2_inv_4 U2313 (.A(n2321), .Y(n2315));
sg13g2_o21ai_1 U2314 (.A1(n4330), .A2(n2319), .B1(n2323), .Y(n2321));
sg13g2_a21oi_2 U2315 (.A1(data_i_93_), .A2(n4308), .B1(n2324), .Y(n2323));
sg13g2_nor2_2 U2316 (.A(n555), .B(n573), .Y(n2324));
sg13g2_inv_4 U2317 (.A(mixcol_data_o_93), .Y(n573));
sg13g2_inv_4 U2318 (.A(subbytes_data_o_93), .Y(n2319));
sg13g2_a21oi_2 U2320 (.A1(n4313), .A2(n2327), .B1(n2328), .Y(n2326));
sg13g2_nor2_2 U2321 (.A(n2329), .B(n4310), .Y(n2328));
sg13g2_o21ai_1 U2322 (.A1(n4167), .A2(n2329), .B1(n2330), .Y(n2327));
sg13g2_a21oi_2 U2323 (.A1(n4315), .A2(n2331), .B1(n2332), .Y(n2330));
sg13g2_nor2_2 U2324 (.A(n4164), .B(n575), .Y(n2332));
sg13g2_inv_4 U2325 (.A(n2331), .Y(n2325));
sg13g2_o21ai_1 U2326 (.A1(n4330), .A2(n2329), .B1(n2333), .Y(n2331));
sg13g2_a21oi_2 U2327 (.A1(data_i_92_), .A2(n4308), .B1(n2334), .Y(n2333));
sg13g2_nor2_2 U2328 (.A(n555), .B(n575), .Y(n2334));
sg13g2_inv_4 U2329 (.A(mixcol_data_o_92), .Y(n575));
sg13g2_inv_4 U2330 (.A(subbytes_data_o_92), .Y(n2329));
sg13g2_a21oi_2 U2332 (.A1(n4313), .A2(n2337), .B1(n2338), .Y(n2336));
sg13g2_nor2_2 U2333 (.A(n2339), .B(n2248), .Y(n2338));
sg13g2_o21ai_1 U2334 (.A1(n4167), .A2(n2339), .B1(n2340), .Y(n2337));
sg13g2_a21oi_2 U2335 (.A1(n4315), .A2(n2341), .B1(n2342), .Y(n2340));
sg13g2_nor2_2 U2336 (.A(n4165), .B(n577), .Y(n2342));
sg13g2_inv_4 U2337 (.A(n2341), .Y(n2335));
sg13g2_o21ai_1 U2338 (.A1(n4330), .A2(n2339), .B1(n2343), .Y(n2341));
sg13g2_a21oi_2 U2339 (.A1(data_i_91_), .A2(n4308), .B1(n2344), .Y(n2343));
sg13g2_nor2_2 U2340 (.A(n555), .B(n577), .Y(n2344));
sg13g2_inv_4 U2341 (.A(mixcol_data_o_91), .Y(n577));
sg13g2_inv_4 U2342 (.A(subbytes_data_o_91), .Y(n2339));
sg13g2_a21oi_2 U2344 (.A1(n4312), .A2(n2347), .B1(n2348), .Y(n2346));
sg13g2_nor2_2 U2345 (.A(n2349), .B(n2248), .Y(n2348));
sg13g2_o21ai_1 U2346 (.A1(n4167), .A2(n2349), .B1(n2350), .Y(n2347));
sg13g2_a21oi_2 U2347 (.A1(n4315), .A2(n2351), .B1(n2352), .Y(n2350));
sg13g2_nor2_2 U2348 (.A(n4165), .B(n579), .Y(n2352));
sg13g2_inv_4 U2349 (.A(n2351), .Y(n2345));
sg13g2_o21ai_1 U2350 (.A1(n4329), .A2(n2349), .B1(n2353), .Y(n2351));
sg13g2_a21oi_2 U2351 (.A1(data_i_90_), .A2(n4308), .B1(n2354), .Y(n2353));
sg13g2_nor2_2 U2352 (.A(n555), .B(n579), .Y(n2354));
sg13g2_inv_4 U2353 (.A(mixcol_data_o_90), .Y(n579));
sg13g2_inv_4 U2354 (.A(subbytes_data_o_90), .Y(n2349));
sg13g2_a21oi_2 U2356 (.A1(n2244), .A2(n2357), .B1(n2358), .Y(n2356));
sg13g2_nor2_2 U2357 (.A(n2359), .B(n2248), .Y(n2358));
sg13g2_o21ai_1 U2358 (.A1(n553), .A2(n2359), .B1(n2360), .Y(n2357));
sg13g2_a21oi_2 U2359 (.A1(n4315), .A2(n2361), .B1(n2362), .Y(n2360));
sg13g2_nor2_2 U2360 (.A(n4165), .B(n581), .Y(n2362));
sg13g2_inv_4 U2361 (.A(n2361), .Y(n2355));
sg13g2_o21ai_1 U2362 (.A1(n4328), .A2(n2359), .B1(n2363), .Y(n2361));
sg13g2_a21oi_2 U2363 (.A1(data_i_8_), .A2(n4308), .B1(n2364), .Y(n2363));
sg13g2_nor2_2 U2364 (.A(n555), .B(n581), .Y(n2364));
sg13g2_inv_4 U2365 (.A(mixcol_data_o_8), .Y(n581));
sg13g2_inv_4 U2366 (.A(subbytes_data_o_8), .Y(n2359));
sg13g2_a21oi_2 U2368 (.A1(n4313), .A2(n2367), .B1(n2368), .Y(n2366));
sg13g2_nor2_2 U2369 (.A(n2369), .B(n4310), .Y(n2368));
sg13g2_o21ai_1 U2370 (.A1(n4167), .A2(n2369), .B1(n2370), .Y(n2367));
sg13g2_a21oi_2 U2371 (.A1(n4315), .A2(n2371), .B1(n2372), .Y(n2370));
sg13g2_nor2_2 U2372 (.A(n4164), .B(n583), .Y(n2372));
sg13g2_inv_4 U2373 (.A(n2371), .Y(n2365));
sg13g2_o21ai_1 U2374 (.A1(n4325), .A2(n2369), .B1(n2373), .Y(n2371));
sg13g2_a21oi_2 U2375 (.A1(data_i_89_), .A2(n4308), .B1(n2374), .Y(n2373));
sg13g2_nor2_2 U2376 (.A(n555), .B(n583), .Y(n2374));
sg13g2_inv_4 U2377 (.A(mixcol_data_o_89), .Y(n583));
sg13g2_inv_4 U2378 (.A(subbytes_data_o_89), .Y(n2369));
sg13g2_a21oi_2 U2380 (.A1(n4313), .A2(n2377), .B1(n2378), .Y(n2376));
sg13g2_nor2_2 U2381 (.A(n2379), .B(n4310), .Y(n2378));
sg13g2_o21ai_1 U2382 (.A1(n553), .A2(n2379), .B1(n2380), .Y(n2377));
sg13g2_a21oi_2 U2383 (.A1(n4315), .A2(n2381), .B1(n2382), .Y(n2380));
sg13g2_nor2_2 U2384 (.A(n4165), .B(n585), .Y(n2382));
sg13g2_inv_4 U2385 (.A(n2381), .Y(n2375));
sg13g2_o21ai_1 U2386 (.A1(n4325), .A2(n2379), .B1(n2383), .Y(n2381));
sg13g2_a21oi_2 U2387 (.A1(data_i_88_), .A2(n4308), .B1(n2384), .Y(n2383));
sg13g2_nor2_2 U2388 (.A(n555), .B(n585), .Y(n2384));
sg13g2_inv_4 U2389 (.A(mixcol_data_o_88), .Y(n585));
sg13g2_inv_4 U2390 (.A(subbytes_data_o_88), .Y(n2379));
sg13g2_a21oi_2 U2392 (.A1(n4313), .A2(n2387), .B1(n2388), .Y(n2386));
sg13g2_nor2_2 U2393 (.A(n2389), .B(n2248), .Y(n2388));
sg13g2_o21ai_1 U2394 (.A1(n553), .A2(n2389), .B1(n2390), .Y(n2387));
sg13g2_a21oi_2 U2395 (.A1(n4315), .A2(n2391), .B1(n2392), .Y(n2390));
sg13g2_nor2_2 U2396 (.A(n4164), .B(n587), .Y(n2392));
sg13g2_inv_4 U2397 (.A(n2391), .Y(n2385));
sg13g2_o21ai_1 U2398 (.A1(n4329), .A2(n2389), .B1(n2393), .Y(n2391));
sg13g2_a21oi_2 U2399 (.A1(data_i_87_), .A2(n4308), .B1(n2394), .Y(n2393));
sg13g2_nor2_2 U2400 (.A(n555), .B(n587), .Y(n2394));
sg13g2_inv_4 U2401 (.A(mixcol_data_o_87), .Y(n587));
sg13g2_inv_4 U2402 (.A(subbytes_data_o_87), .Y(n2389));
sg13g2_a21oi_2 U2404 (.A1(n2244), .A2(n2397), .B1(n2398), .Y(n2396));
sg13g2_nor2_2 U2405 (.A(n2399), .B(n2248), .Y(n2398));
sg13g2_o21ai_1 U2406 (.A1(n4167), .A2(n2399), .B1(n2400), .Y(n2397));
sg13g2_a21oi_2 U2407 (.A1(n4315), .A2(n2401), .B1(n2402), .Y(n2400));
sg13g2_nor2_2 U2408 (.A(n4165), .B(n589), .Y(n2402));
sg13g2_inv_4 U2409 (.A(n2401), .Y(n2395));
sg13g2_o21ai_1 U2410 (.A1(n4325), .A2(n2399), .B1(n2403), .Y(n2401));
sg13g2_a21oi_2 U2411 (.A1(data_i_86_), .A2(n4308), .B1(n2404), .Y(n2403));
sg13g2_nor2_2 U2412 (.A(n555), .B(n589), .Y(n2404));
sg13g2_inv_4 U2413 (.A(mixcol_data_o_86), .Y(n589));
sg13g2_inv_4 U2414 (.A(subbytes_data_o_86), .Y(n2399));
sg13g2_a21oi_2 U2416 (.A1(n4313), .A2(n2407), .B1(n2408), .Y(n2406));
sg13g2_nor2_2 U2417 (.A(n2409), .B(n4310), .Y(n2408));
sg13g2_o21ai_1 U2418 (.A1(n4167), .A2(n2409), .B1(n2410), .Y(n2407));
sg13g2_a21oi_2 U2419 (.A1(n4315), .A2(n2411), .B1(n2412), .Y(n2410));
sg13g2_nor2_2 U2420 (.A(n4164), .B(n591), .Y(n2412));
sg13g2_inv_4 U2421 (.A(n2411), .Y(n2405));
sg13g2_o21ai_1 U2422 (.A1(n4330), .A2(n2409), .B1(n2413), .Y(n2411));
sg13g2_a21oi_2 U2423 (.A1(data_i_85_), .A2(n4308), .B1(n2414), .Y(n2413));
sg13g2_nor2_2 U2424 (.A(n555), .B(n591), .Y(n2414));
sg13g2_inv_4 U2425 (.A(mixcol_data_o_85), .Y(n591));
sg13g2_inv_4 U2426 (.A(subbytes_data_o_85), .Y(n2409));
sg13g2_a21oi_2 U2428 (.A1(n4313), .A2(n2417), .B1(n2418), .Y(n2416));
sg13g2_nor2_2 U2429 (.A(n2419), .B(n2248), .Y(n2418));
sg13g2_o21ai_1 U2430 (.A1(n553), .A2(n2419), .B1(n2420), .Y(n2417));
sg13g2_a21oi_2 U2431 (.A1(n4315), .A2(n2421), .B1(n2422), .Y(n2420));
sg13g2_nor2_2 U2432 (.A(n4164), .B(n593), .Y(n2422));
sg13g2_inv_4 U2433 (.A(n2421), .Y(n2415));
sg13g2_o21ai_1 U2434 (.A1(n4327), .A2(n2419), .B1(n2423), .Y(n2421));
sg13g2_a21oi_2 U2435 (.A1(data_i_84_), .A2(n4308), .B1(n2424), .Y(n2423));
sg13g2_nor2_2 U2436 (.A(n555), .B(n593), .Y(n2424));
sg13g2_inv_4 U2437 (.A(mixcol_data_o_84), .Y(n593));
sg13g2_inv_4 U2438 (.A(subbytes_data_o_84), .Y(n2419));
sg13g2_a21oi_2 U2440 (.A1(n4313), .A2(n2427), .B1(n2428), .Y(n2426));
sg13g2_nor2_2 U2441 (.A(n2429), .B(n4310), .Y(n2428));
sg13g2_o21ai_1 U2442 (.A1(n553), .A2(n2429), .B1(n2430), .Y(n2427));
sg13g2_a21oi_2 U2443 (.A1(n4315), .A2(n2431), .B1(n2432), .Y(n2430));
sg13g2_nor2_2 U2444 (.A(n4165), .B(n595), .Y(n2432));
sg13g2_inv_4 U2445 (.A(n2431), .Y(n2425));
sg13g2_o21ai_1 U2446 (.A1(n4326), .A2(n2429), .B1(n2433), .Y(n2431));
sg13g2_a21oi_2 U2447 (.A1(data_i_83_), .A2(n4308), .B1(n2434), .Y(n2433));
sg13g2_nor2_2 U2448 (.A(n555), .B(n595), .Y(n2434));
sg13g2_inv_4 U2449 (.A(mixcol_data_o_83), .Y(n595));
sg13g2_inv_4 U2450 (.A(subbytes_data_o_83), .Y(n2429));
sg13g2_a21oi_2 U2452 (.A1(n4313), .A2(n2437), .B1(n2438), .Y(n2436));
sg13g2_nor2_2 U2453 (.A(n2439), .B(n4310), .Y(n2438));
sg13g2_o21ai_1 U2454 (.A1(n4167), .A2(n2439), .B1(n2440), .Y(n2437));
sg13g2_a21oi_2 U2455 (.A1(n4315), .A2(n2441), .B1(n2442), .Y(n2440));
sg13g2_nor2_2 U2456 (.A(n4165), .B(n597), .Y(n2442));
sg13g2_inv_4 U2457 (.A(n2441), .Y(n2435));
sg13g2_o21ai_1 U2458 (.A1(n4326), .A2(n2439), .B1(n2443), .Y(n2441));
sg13g2_a21oi_2 U2459 (.A1(data_i_82_), .A2(n4308), .B1(n2444), .Y(n2443));
sg13g2_nor2_2 U2460 (.A(n555), .B(n597), .Y(n2444));
sg13g2_inv_4 U2461 (.A(mixcol_data_o_82), .Y(n597));
sg13g2_inv_4 U2462 (.A(subbytes_data_o_82), .Y(n2439));
sg13g2_a21oi_2 U2464 (.A1(n4313), .A2(n2447), .B1(n2448), .Y(n2446));
sg13g2_nor2_2 U2465 (.A(n2449), .B(n2248), .Y(n2448));
sg13g2_o21ai_1 U2466 (.A1(n4167), .A2(n2449), .B1(n2450), .Y(n2447));
sg13g2_a21oi_2 U2467 (.A1(n4315), .A2(n2451), .B1(n2452), .Y(n2450));
sg13g2_nor2_2 U2468 (.A(n4165), .B(n599), .Y(n2452));
sg13g2_inv_4 U2469 (.A(n2451), .Y(n2445));
sg13g2_o21ai_1 U2470 (.A1(n4325), .A2(n2449), .B1(n2453), .Y(n2451));
sg13g2_a21oi_2 U2471 (.A1(data_i_81_), .A2(n4307), .B1(n2454), .Y(n2453));
sg13g2_nor2_2 U2472 (.A(n555), .B(n599), .Y(n2454));
sg13g2_inv_4 U2473 (.A(mixcol_data_o_81), .Y(n599));
sg13g2_inv_4 U2474 (.A(subbytes_data_o_81), .Y(n2449));
sg13g2_a21oi_2 U2476 (.A1(n4313), .A2(n2457), .B1(n2458), .Y(n2456));
sg13g2_nor2_2 U2477 (.A(n2459), .B(n4310), .Y(n2458));
sg13g2_o21ai_1 U2478 (.A1(n553), .A2(n2459), .B1(n2460), .Y(n2457));
sg13g2_a21oi_2 U2479 (.A1(n4315), .A2(n2461), .B1(n2462), .Y(n2460));
sg13g2_nor2_2 U2480 (.A(n4164), .B(n601), .Y(n2462));
sg13g2_inv_4 U2481 (.A(n2461), .Y(n2455));
sg13g2_o21ai_1 U2482 (.A1(n4330), .A2(n2459), .B1(n2463), .Y(n2461));
sg13g2_a21oi_2 U2483 (.A1(data_i_80_), .A2(n4308), .B1(n2464), .Y(n2463));
sg13g2_nor2_2 U2484 (.A(n555), .B(n601), .Y(n2464));
sg13g2_inv_4 U2485 (.A(mixcol_data_o_80), .Y(n601));
sg13g2_inv_4 U2486 (.A(subbytes_data_o_80), .Y(n2459));
sg13g2_a21oi_2 U2488 (.A1(n4313), .A2(n2467), .B1(n2468), .Y(n2466));
sg13g2_nor2_2 U2489 (.A(n2469), .B(n2248), .Y(n2468));
sg13g2_o21ai_1 U2490 (.A1(n4167), .A2(n2469), .B1(n2470), .Y(n2467));
sg13g2_a21oi_2 U2491 (.A1(n4315), .A2(n2471), .B1(n2472), .Y(n2470));
sg13g2_nor2_2 U2492 (.A(n4164), .B(n603), .Y(n2472));
sg13g2_inv_4 U2493 (.A(n2471), .Y(n2465));
sg13g2_o21ai_1 U2494 (.A1(n4329), .A2(n2469), .B1(n2473), .Y(n2471));
sg13g2_a21oi_2 U2495 (.A1(data_i_7_), .A2(n4307), .B1(n2474), .Y(n2473));
sg13g2_nor2_2 U2496 (.A(n555), .B(n603), .Y(n2474));
sg13g2_inv_4 U2497 (.A(mixcol_data_o_7), .Y(n603));
sg13g2_inv_4 U2498 (.A(subbytes_data_o_7), .Y(n2469));
sg13g2_a21oi_2 U2500 (.A1(n4313), .A2(n2477), .B1(n2478), .Y(n2476));
sg13g2_nor2_2 U2501 (.A(n2479), .B(n2248), .Y(n2478));
sg13g2_o21ai_1 U2502 (.A1(n553), .A2(n2479), .B1(n2480), .Y(n2477));
sg13g2_a21oi_2 U2503 (.A1(n4315), .A2(n2481), .B1(n2482), .Y(n2480));
sg13g2_nor2_2 U2504 (.A(n4165), .B(n605), .Y(n2482));
sg13g2_inv_4 U2505 (.A(n2481), .Y(n2475));
sg13g2_o21ai_1 U2506 (.A1(n4328), .A2(n2479), .B1(n2483), .Y(n2481));
sg13g2_a21oi_2 U2507 (.A1(data_i_79_), .A2(n4308), .B1(n2484), .Y(n2483));
sg13g2_nor2_2 U2508 (.A(n555), .B(n605), .Y(n2484));
sg13g2_inv_4 U2509 (.A(mixcol_data_o_79), .Y(n605));
sg13g2_inv_4 U2510 (.A(subbytes_data_o_79), .Y(n2479));
sg13g2_a21oi_2 U2512 (.A1(n4313), .A2(n2487), .B1(n2488), .Y(n2486));
sg13g2_nor2_2 U2513 (.A(n2489), .B(n4310), .Y(n2488));
sg13g2_o21ai_1 U2514 (.A1(n4167), .A2(n2489), .B1(n2490), .Y(n2487));
sg13g2_a21oi_2 U2515 (.A1(n4315), .A2(n2491), .B1(n2492), .Y(n2490));
sg13g2_nor2_2 U2516 (.A(n4164), .B(n607), .Y(n2492));
sg13g2_inv_4 U2517 (.A(n2491), .Y(n2485));
sg13g2_o21ai_1 U2518 (.A1(n4325), .A2(n2489), .B1(n2493), .Y(n2491));
sg13g2_a21oi_2 U2519 (.A1(data_i_78_), .A2(n4308), .B1(n2494), .Y(n2493));
sg13g2_nor2_2 U2520 (.A(n555), .B(n607), .Y(n2494));
sg13g2_inv_4 U2521 (.A(mixcol_data_o_78), .Y(n607));
sg13g2_inv_4 U2522 (.A(subbytes_data_o_78), .Y(n2489));
sg13g2_a21oi_2 U2524 (.A1(n4313), .A2(n2497), .B1(n2498), .Y(n2496));
sg13g2_nor2_2 U2525 (.A(n2499), .B(n2248), .Y(n2498));
sg13g2_o21ai_1 U2526 (.A1(n4167), .A2(n2499), .B1(n2500), .Y(n2497));
sg13g2_a21oi_2 U2527 (.A1(n4315), .A2(n2501), .B1(n2502), .Y(n2500));
sg13g2_nor2_2 U2528 (.A(n4165), .B(n609), .Y(n2502));
sg13g2_inv_4 U2529 (.A(n2501), .Y(n2495));
sg13g2_o21ai_1 U2530 (.A1(n4327), .A2(n2499), .B1(n2503), .Y(n2501));
sg13g2_a21oi_2 U2531 (.A1(data_i_77_), .A2(n4308), .B1(n2504), .Y(n2503));
sg13g2_nor2_2 U2532 (.A(n555), .B(n609), .Y(n2504));
sg13g2_inv_4 U2533 (.A(mixcol_data_o_77), .Y(n609));
sg13g2_inv_4 U2534 (.A(subbytes_data_o_77), .Y(n2499));
sg13g2_a21oi_2 U2536 (.A1(n4313), .A2(n2507), .B1(n2508), .Y(n2506));
sg13g2_nor2_2 U2537 (.A(n2509), .B(n2248), .Y(n2508));
sg13g2_o21ai_1 U2538 (.A1(n553), .A2(n2509), .B1(n2510), .Y(n2507));
sg13g2_a21oi_2 U2539 (.A1(n4315), .A2(n2511), .B1(n2512), .Y(n2510));
sg13g2_nor2_2 U2540 (.A(n4164), .B(n611), .Y(n2512));
sg13g2_inv_4 U2541 (.A(n2511), .Y(n2505));
sg13g2_o21ai_1 U2542 (.A1(n4328), .A2(n2509), .B1(n2513), .Y(n2511));
sg13g2_a21oi_2 U2543 (.A1(data_i_76_), .A2(n4307), .B1(n2514), .Y(n2513));
sg13g2_nor2_2 U2544 (.A(n555), .B(n611), .Y(n2514));
sg13g2_inv_4 U2545 (.A(mixcol_data_o_76), .Y(n611));
sg13g2_inv_4 U2546 (.A(subbytes_data_o_76), .Y(n2509));
sg13g2_a21oi_2 U2548 (.A1(n4313), .A2(n2517), .B1(n2518), .Y(n2516));
sg13g2_nor2_2 U2549 (.A(n2519), .B(n2248), .Y(n2518));
sg13g2_o21ai_1 U2550 (.A1(n553), .A2(n2519), .B1(n2520), .Y(n2517));
sg13g2_a21oi_2 U2551 (.A1(n4315), .A2(n2521), .B1(n2522), .Y(n2520));
sg13g2_nor2_2 U2552 (.A(n4165), .B(n613), .Y(n2522));
sg13g2_inv_4 U2553 (.A(n2521), .Y(n2515));
sg13g2_o21ai_1 U2554 (.A1(n4329), .A2(n2519), .B1(n2523), .Y(n2521));
sg13g2_a21oi_2 U2555 (.A1(data_i_75_), .A2(n4308), .B1(n2524), .Y(n2523));
sg13g2_nor2_2 U2556 (.A(n555), .B(n613), .Y(n2524));
sg13g2_inv_4 U2557 (.A(mixcol_data_o_75), .Y(n613));
sg13g2_inv_4 U2558 (.A(subbytes_data_o_75), .Y(n2519));
sg13g2_a21oi_2 U2560 (.A1(n2244), .A2(n2527), .B1(n2528), .Y(n2526));
sg13g2_nor2_2 U2561 (.A(n2529), .B(n2248), .Y(n2528));
sg13g2_o21ai_1 U2562 (.A1(n4167), .A2(n2529), .B1(n2530), .Y(n2527));
sg13g2_a21oi_2 U2563 (.A1(n4315), .A2(n2531), .B1(n2532), .Y(n2530));
sg13g2_nor2_2 U2564 (.A(n4164), .B(n615), .Y(n2532));
sg13g2_inv_4 U2565 (.A(n2531), .Y(n2525));
sg13g2_o21ai_1 U2566 (.A1(n4325), .A2(n2529), .B1(n2533), .Y(n2531));
sg13g2_a21oi_2 U2567 (.A1(data_i_74_), .A2(n4307), .B1(n2534), .Y(n2533));
sg13g2_nor2_2 U2568 (.A(n555), .B(n615), .Y(n2534));
sg13g2_inv_4 U2569 (.A(mixcol_data_o_74), .Y(n615));
sg13g2_inv_4 U2570 (.A(subbytes_data_o_74), .Y(n2529));
sg13g2_o21ai_1 U2571 (.A1(state), .A2(n2535), .B1(n2536), .Y(addroundkey_data_i_73));
sg13g2_a21oi_2 U2572 (.A1(n2244), .A2(n2537), .B1(n2538), .Y(n2536));
sg13g2_nor2_2 U2573 (.A(n2539), .B(n4310), .Y(n2538));
sg13g2_o21ai_1 U2574 (.A1(n553), .A2(n2539), .B1(n2540), .Y(n2537));
sg13g2_a21oi_2 U2575 (.A1(n4315), .A2(n2541), .B1(n2542), .Y(n2540));
sg13g2_nor2_2 U2576 (.A(n4164), .B(n617), .Y(n2542));
sg13g2_inv_4 U2577 (.A(n2541), .Y(n2535));
sg13g2_o21ai_1 U2578 (.A1(n4326), .A2(n2539), .B1(n2543), .Y(n2541));
sg13g2_a21oi_2 U2579 (.A1(data_i_73_), .A2(n4308), .B1(n2544), .Y(n2543));
sg13g2_nor2_2 U2580 (.A(n555), .B(n617), .Y(n2544));
sg13g2_inv_4 U2581 (.A(mixcol_data_o_73), .Y(n617));
sg13g2_inv_4 U2582 (.A(subbytes_data_o_73), .Y(n2539));
sg13g2_a21oi_2 U2584 (.A1(n2244), .A2(n2547), .B1(n2548), .Y(n2546));
sg13g2_nor2_2 U2585 (.A(n2549), .B(n2248), .Y(n2548));
sg13g2_o21ai_1 U2586 (.A1(n4167), .A2(n2549), .B1(n2550), .Y(n2547));
sg13g2_a21oi_2 U2587 (.A1(n4315), .A2(n2551), .B1(n2552), .Y(n2550));
sg13g2_nor2_2 U2588 (.A(n4164), .B(n619), .Y(n2552));
sg13g2_inv_4 U2589 (.A(n2551), .Y(n2545));
sg13g2_o21ai_1 U2590 (.A1(n4327), .A2(n2549), .B1(n2553), .Y(n2551));
sg13g2_a21oi_2 U2591 (.A1(data_i_72_), .A2(n4307), .B1(n2554), .Y(n2553));
sg13g2_nor2_2 U2592 (.A(n555), .B(n619), .Y(n2554));
sg13g2_inv_4 U2593 (.A(mixcol_data_o_72), .Y(n619));
sg13g2_inv_4 U2594 (.A(subbytes_data_o_72), .Y(n2549));
sg13g2_a21oi_2 U2596 (.A1(n2244), .A2(n2557), .B1(n2558), .Y(n2556));
sg13g2_nor2_2 U2597 (.A(n2559), .B(n2248), .Y(n2558));
sg13g2_o21ai_1 U2598 (.A1(n4167), .A2(n2559), .B1(n2560), .Y(n2557));
sg13g2_a21oi_2 U2599 (.A1(n4315), .A2(n2561), .B1(n2562), .Y(n2560));
sg13g2_nor2_2 U2600 (.A(n4165), .B(n621), .Y(n2562));
sg13g2_inv_4 U2601 (.A(n2561), .Y(n2555));
sg13g2_o21ai_1 U2602 (.A1(n4330), .A2(n2559), .B1(n2563), .Y(n2561));
sg13g2_a21oi_2 U2603 (.A1(data_i_71_), .A2(n4307), .B1(n2564), .Y(n2563));
sg13g2_nor2_2 U2604 (.A(n555), .B(n621), .Y(n2564));
sg13g2_inv_4 U2605 (.A(mixcol_data_o_71), .Y(n621));
sg13g2_inv_4 U2606 (.A(subbytes_data_o_71), .Y(n2559));
sg13g2_a21oi_2 U2608 (.A1(n4312), .A2(n2567), .B1(n2568), .Y(n2566));
sg13g2_nor2_2 U2609 (.A(n2569), .B(n2248), .Y(n2568));
sg13g2_o21ai_1 U2610 (.A1(n553), .A2(n2569), .B1(n2570), .Y(n2567));
sg13g2_a21oi_2 U2611 (.A1(n4315), .A2(n2571), .B1(n2572), .Y(n2570));
sg13g2_nor2_2 U2612 (.A(n4164), .B(n623), .Y(n2572));
sg13g2_inv_4 U2613 (.A(n2571), .Y(n2565));
sg13g2_o21ai_1 U2614 (.A1(n4327), .A2(n2569), .B1(n2573), .Y(n2571));
sg13g2_a21oi_2 U2615 (.A1(data_i_70_), .A2(n4308), .B1(n2574), .Y(n2573));
sg13g2_nor2_2 U2616 (.A(n555), .B(n623), .Y(n2574));
sg13g2_inv_4 U2617 (.A(mixcol_data_o_70), .Y(n623));
sg13g2_inv_4 U2618 (.A(subbytes_data_o_70), .Y(n2569));
sg13g2_a21oi_2 U2620 (.A1(n2244), .A2(n2577), .B1(n2578), .Y(n2576));
sg13g2_nor2_2 U2621 (.A(n2579), .B(n2248), .Y(n2578));
sg13g2_o21ai_1 U2622 (.A1(n553), .A2(n2579), .B1(n2580), .Y(n2577));
sg13g2_a21oi_2 U2623 (.A1(n4315), .A2(n2581), .B1(n2582), .Y(n2580));
sg13g2_nor2_2 U2624 (.A(n4165), .B(n625), .Y(n2582));
sg13g2_inv_4 U2625 (.A(n2581), .Y(n2575));
sg13g2_o21ai_1 U2626 (.A1(n4329), .A2(n2579), .B1(n2583), .Y(n2581));
sg13g2_a21oi_2 U2627 (.A1(data_i_6_), .A2(n4307), .B1(n2584), .Y(n2583));
sg13g2_nor2_2 U2628 (.A(n555), .B(n625), .Y(n2584));
sg13g2_inv_4 U2629 (.A(mixcol_data_o_6), .Y(n625));
sg13g2_inv_4 U2630 (.A(subbytes_data_o_6), .Y(n2579));
sg13g2_o21ai_1 U2631 (.A1(state), .A2(n2585), .B1(n2586), .Y(addroundkey_data_i_69));
sg13g2_a21oi_2 U2632 (.A1(n4313), .A2(n2587), .B1(n2588), .Y(n2586));
sg13g2_nor2_2 U2633 (.A(n2589), .B(n4310), .Y(n2588));
sg13g2_o21ai_1 U2634 (.A1(n553), .A2(n2589), .B1(n2590), .Y(n2587));
sg13g2_a21oi_2 U2635 (.A1(n4315), .A2(n2591), .B1(n2592), .Y(n2590));
sg13g2_nor2_2 U2636 (.A(n4165), .B(n627), .Y(n2592));
sg13g2_inv_4 U2637 (.A(n2591), .Y(n2585));
sg13g2_o21ai_1 U2638 (.A1(n4326), .A2(n2589), .B1(n2593), .Y(n2591));
sg13g2_a21oi_2 U2639 (.A1(data_i_69_), .A2(n4308), .B1(n2594), .Y(n2593));
sg13g2_nor2_2 U2640 (.A(n555), .B(n627), .Y(n2594));
sg13g2_inv_4 U2641 (.A(mixcol_data_o_69), .Y(n627));
sg13g2_inv_4 U2642 (.A(subbytes_data_o_69), .Y(n2589));
sg13g2_a21oi_2 U2644 (.A1(n4313), .A2(n2597), .B1(n2598), .Y(n2596));
sg13g2_nor2_2 U2645 (.A(n2599), .B(n4310), .Y(n2598));
sg13g2_o21ai_1 U2646 (.A1(n553), .A2(n2599), .B1(n2600), .Y(n2597));
sg13g2_a21oi_2 U2647 (.A1(n4315), .A2(n2601), .B1(n2602), .Y(n2600));
sg13g2_nor2_2 U2648 (.A(n4164), .B(n629), .Y(n2602));
sg13g2_inv_4 U2649 (.A(n2601), .Y(n2595));
sg13g2_o21ai_1 U2650 (.A1(n4327), .A2(n2599), .B1(n2603), .Y(n2601));
sg13g2_a21oi_2 U2651 (.A1(data_i_68_), .A2(n4308), .B1(n2604), .Y(n2603));
sg13g2_nor2_2 U2652 (.A(n555), .B(n629), .Y(n2604));
sg13g2_inv_4 U2653 (.A(mixcol_data_o_68), .Y(n629));
sg13g2_inv_4 U2654 (.A(subbytes_data_o_68), .Y(n2599));
sg13g2_a21oi_2 U2656 (.A1(n4312), .A2(n2607), .B1(n2608), .Y(n2606));
sg13g2_nor2_2 U2657 (.A(n2609), .B(n4310), .Y(n2608));
sg13g2_o21ai_1 U2658 (.A1(n553), .A2(n2609), .B1(n2610), .Y(n2607));
sg13g2_a21oi_2 U2659 (.A1(n4315), .A2(n2611), .B1(n2612), .Y(n2610));
sg13g2_nor2_2 U2660 (.A(n4164), .B(n631), .Y(n2612));
sg13g2_inv_4 U2661 (.A(n2611), .Y(n2605));
sg13g2_o21ai_1 U2662 (.A1(n4328), .A2(n2609), .B1(n2613), .Y(n2611));
sg13g2_a21oi_2 U2663 (.A1(data_i_67_), .A2(n4308), .B1(n2614), .Y(n2613));
sg13g2_nor2_2 U2664 (.A(n555), .B(n631), .Y(n2614));
sg13g2_inv_4 U2665 (.A(mixcol_data_o_67), .Y(n631));
sg13g2_inv_4 U2666 (.A(subbytes_data_o_67), .Y(n2609));
sg13g2_a21oi_2 U2668 (.A1(n4313), .A2(n2617), .B1(n2618), .Y(n2616));
sg13g2_nor2_2 U2669 (.A(n2619), .B(n4310), .Y(n2618));
sg13g2_o21ai_1 U2670 (.A1(n553), .A2(n2619), .B1(n2620), .Y(n2617));
sg13g2_a21oi_2 U2671 (.A1(n4315), .A2(n2621), .B1(n2622), .Y(n2620));
sg13g2_nor2_2 U2672 (.A(n4165), .B(n633), .Y(n2622));
sg13g2_inv_4 U2673 (.A(n2621), .Y(n2615));
sg13g2_o21ai_1 U2674 (.A1(n4326), .A2(n2619), .B1(n2623), .Y(n2621));
sg13g2_a21oi_2 U2675 (.A1(data_i_66_), .A2(n4307), .B1(n2624), .Y(n2623));
sg13g2_nor2_2 U2676 (.A(n555), .B(n633), .Y(n2624));
sg13g2_inv_4 U2677 (.A(mixcol_data_o_66), .Y(n633));
sg13g2_inv_4 U2678 (.A(subbytes_data_o_66), .Y(n2619));
sg13g2_a21oi_2 U2680 (.A1(n4312), .A2(n2627), .B1(n2628), .Y(n2626));
sg13g2_nor2_2 U2681 (.A(n2629), .B(n4310), .Y(n2628));
sg13g2_o21ai_1 U2682 (.A1(n4167), .A2(n2629), .B1(n2630), .Y(n2627));
sg13g2_a21oi_2 U2683 (.A1(n4315), .A2(n2631), .B1(n2632), .Y(n2630));
sg13g2_nor2_2 U2684 (.A(n4165), .B(n635), .Y(n2632));
sg13g2_inv_4 U2685 (.A(n2631), .Y(n2625));
sg13g2_o21ai_1 U2686 (.A1(n4327), .A2(n2629), .B1(n2633), .Y(n2631));
sg13g2_a21oi_2 U2687 (.A1(data_i_65_), .A2(n4308), .B1(n2634), .Y(n2633));
sg13g2_nor2_2 U2688 (.A(n555), .B(n635), .Y(n2634));
sg13g2_inv_4 U2689 (.A(mixcol_data_o_65), .Y(n635));
sg13g2_inv_4 U2690 (.A(subbytes_data_o_65), .Y(n2629));
sg13g2_a21oi_2 U2692 (.A1(n4313), .A2(n2637), .B1(n2638), .Y(n2636));
sg13g2_nor2_2 U2693 (.A(n2639), .B(n2248), .Y(n2638));
sg13g2_o21ai_1 U2694 (.A1(n4167), .A2(n2639), .B1(n2640), .Y(n2637));
sg13g2_a21oi_2 U2695 (.A1(n4315), .A2(n2641), .B1(n2642), .Y(n2640));
sg13g2_nor2_2 U2696 (.A(n4165), .B(n637), .Y(n2642));
sg13g2_inv_4 U2697 (.A(n2641), .Y(n2635));
sg13g2_o21ai_1 U2698 (.A1(n4330), .A2(n2639), .B1(n2643), .Y(n2641));
sg13g2_a21oi_2 U2699 (.A1(data_i_64_), .A2(n4308), .B1(n2644), .Y(n2643));
sg13g2_nor2_2 U2700 (.A(n555), .B(n637), .Y(n2644));
sg13g2_inv_4 U2701 (.A(mixcol_data_o_64), .Y(n637));
sg13g2_inv_4 U2702 (.A(subbytes_data_o_64), .Y(n2639));
sg13g2_a21oi_2 U2704 (.A1(n4313), .A2(n2647), .B1(n2648), .Y(n2646));
sg13g2_nor2_2 U2705 (.A(n2649), .B(n4310), .Y(n2648));
sg13g2_o21ai_1 U2706 (.A1(n4167), .A2(n2649), .B1(n2650), .Y(n2647));
sg13g2_a21oi_2 U2707 (.A1(n4315), .A2(n2651), .B1(n2652), .Y(n2650));
sg13g2_nor2_2 U2708 (.A(n4165), .B(n639), .Y(n2652));
sg13g2_inv_4 U2709 (.A(n2651), .Y(n2645));
sg13g2_o21ai_1 U2710 (.A1(n4327), .A2(n2649), .B1(n2653), .Y(n2651));
sg13g2_a21oi_2 U2711 (.A1(data_i_63_), .A2(n4308), .B1(n2654), .Y(n2653));
sg13g2_nor2_2 U2712 (.A(n555), .B(n639), .Y(n2654));
sg13g2_inv_4 U2713 (.A(mixcol_data_o_63), .Y(n639));
sg13g2_inv_4 U2714 (.A(subbytes_data_o_63), .Y(n2649));
sg13g2_a21oi_2 U2716 (.A1(n4313), .A2(n2657), .B1(n2658), .Y(n2656));
sg13g2_nor2_2 U2717 (.A(n2659), .B(n4310), .Y(n2658));
sg13g2_o21ai_1 U2718 (.A1(n553), .A2(n2659), .B1(n2660), .Y(n2657));
sg13g2_a21oi_2 U2719 (.A1(n4315), .A2(n2661), .B1(n2662), .Y(n2660));
sg13g2_nor2_2 U2720 (.A(n4165), .B(n641), .Y(n2662));
sg13g2_inv_4 U2721 (.A(n2661), .Y(n2655));
sg13g2_o21ai_1 U2722 (.A1(n4328), .A2(n2659), .B1(n2663), .Y(n2661));
sg13g2_a21oi_2 U2723 (.A1(data_i_62_), .A2(n4308), .B1(n2664), .Y(n2663));
sg13g2_nor2_2 U2724 (.A(n555), .B(n641), .Y(n2664));
sg13g2_inv_4 U2725 (.A(mixcol_data_o_62), .Y(n641));
sg13g2_inv_4 U2726 (.A(subbytes_data_o_62), .Y(n2659));
sg13g2_a21oi_2 U2728 (.A1(n4313), .A2(n2667), .B1(n2668), .Y(n2666));
sg13g2_nor2_2 U2729 (.A(n2669), .B(n4310), .Y(n2668));
sg13g2_o21ai_1 U2730 (.A1(n4167), .A2(n2669), .B1(n2670), .Y(n2667));
sg13g2_a21oi_2 U2731 (.A1(n4315), .A2(n2671), .B1(n2672), .Y(n2670));
sg13g2_nor2_2 U2732 (.A(n4164), .B(n643), .Y(n2672));
sg13g2_inv_4 U2733 (.A(n2671), .Y(n2665));
sg13g2_o21ai_1 U2734 (.A1(n4329), .A2(n2669), .B1(n2673), .Y(n2671));
sg13g2_a21oi_2 U2735 (.A1(data_i_61_), .A2(n4308), .B1(n2674), .Y(n2673));
sg13g2_nor2_2 U2736 (.A(n555), .B(n643), .Y(n2674));
sg13g2_inv_4 U2737 (.A(mixcol_data_o_61), .Y(n643));
sg13g2_inv_4 U2738 (.A(subbytes_data_o_61), .Y(n2669));
sg13g2_a21oi_2 U2740 (.A1(n4312), .A2(n2677), .B1(n2678), .Y(n2676));
sg13g2_nor2_2 U2741 (.A(n2679), .B(n4310), .Y(n2678));
sg13g2_o21ai_1 U2742 (.A1(n553), .A2(n2679), .B1(n2680), .Y(n2677));
sg13g2_a21oi_2 U2743 (.A1(n4315), .A2(n2681), .B1(n2682), .Y(n2680));
sg13g2_nor2_2 U2744 (.A(n4165), .B(n645), .Y(n2682));
sg13g2_inv_4 U2745 (.A(n2681), .Y(n2675));
sg13g2_o21ai_1 U2746 (.A1(n4328), .A2(n2679), .B1(n2683), .Y(n2681));
sg13g2_a21oi_2 U2747 (.A1(data_i_60_), .A2(n4308), .B1(n2684), .Y(n2683));
sg13g2_nor2_2 U2748 (.A(n555), .B(n645), .Y(n2684));
sg13g2_inv_4 U2749 (.A(mixcol_data_o_60), .Y(n645));
sg13g2_inv_4 U2750 (.A(subbytes_data_o_60), .Y(n2679));
sg13g2_a21oi_2 U2752 (.A1(n4312), .A2(n2687), .B1(n2688), .Y(n2686));
sg13g2_nor2_2 U2753 (.A(n2689), .B(n4310), .Y(n2688));
sg13g2_o21ai_1 U2754 (.A1(n553), .A2(n2689), .B1(n2690), .Y(n2687));
sg13g2_a21oi_2 U2755 (.A1(n4315), .A2(n2691), .B1(n2692), .Y(n2690));
sg13g2_nor2_2 U2756 (.A(n4165), .B(n647), .Y(n2692));
sg13g2_inv_4 U2757 (.A(n2691), .Y(n2685));
sg13g2_o21ai_1 U2758 (.A1(n4330), .A2(n2689), .B1(n2693), .Y(n2691));
sg13g2_a21oi_2 U2759 (.A1(data_i_5_), .A2(n4308), .B1(n2694), .Y(n2693));
sg13g2_nor2_2 U2760 (.A(n555), .B(n647), .Y(n2694));
sg13g2_inv_4 U2761 (.A(mixcol_data_o_5), .Y(n647));
sg13g2_inv_4 U2762 (.A(subbytes_data_o_5), .Y(n2689));
sg13g2_a21oi_2 U2764 (.A1(n4313), .A2(n2697), .B1(n2698), .Y(n2696));
sg13g2_nor2_2 U2765 (.A(n2699), .B(n2248), .Y(n2698));
sg13g2_o21ai_1 U2766 (.A1(n553), .A2(n2699), .B1(n2700), .Y(n2697));
sg13g2_a21oi_2 U2767 (.A1(n4315), .A2(n2701), .B1(n2702), .Y(n2700));
sg13g2_nor2_2 U2768 (.A(n4164), .B(n649), .Y(n2702));
sg13g2_inv_4 U2769 (.A(n2701), .Y(n2695));
sg13g2_o21ai_1 U2770 (.A1(n4329), .A2(n2699), .B1(n2703), .Y(n2701));
sg13g2_a21oi_2 U2771 (.A1(data_i_59_), .A2(n4308), .B1(n2704), .Y(n2703));
sg13g2_nor2_2 U2772 (.A(n555), .B(n649), .Y(n2704));
sg13g2_inv_4 U2773 (.A(mixcol_data_o_59), .Y(n649));
sg13g2_inv_4 U2774 (.A(subbytes_data_o_59), .Y(n2699));
sg13g2_a21oi_2 U2776 (.A1(n4313), .A2(n2707), .B1(n2708), .Y(n2706));
sg13g2_nor2_2 U2777 (.A(n2709), .B(n4310), .Y(n2708));
sg13g2_o21ai_1 U2778 (.A1(n4167), .A2(n2709), .B1(n2710), .Y(n2707));
sg13g2_a21oi_2 U2779 (.A1(n4315), .A2(n2711), .B1(n2712), .Y(n2710));
sg13g2_nor2_2 U2780 (.A(n4165), .B(n651), .Y(n2712));
sg13g2_inv_4 U2781 (.A(n2711), .Y(n2705));
sg13g2_o21ai_1 U2782 (.A1(n4327), .A2(n2709), .B1(n2713), .Y(n2711));
sg13g2_a21oi_2 U2783 (.A1(data_i_58_), .A2(n4308), .B1(n2714), .Y(n2713));
sg13g2_nor2_2 U2784 (.A(n555), .B(n651), .Y(n2714));
sg13g2_inv_4 U2785 (.A(mixcol_data_o_58), .Y(n651));
sg13g2_inv_4 U2786 (.A(subbytes_data_o_58), .Y(n2709));
sg13g2_a21oi_2 U2788 (.A1(n4313), .A2(n2717), .B1(n2718), .Y(n2716));
sg13g2_nor2_2 U2789 (.A(n2719), .B(n2248), .Y(n2718));
sg13g2_o21ai_1 U2790 (.A1(n553), .A2(n2719), .B1(n2720), .Y(n2717));
sg13g2_a21oi_2 U2791 (.A1(n4315), .A2(n2721), .B1(n2722), .Y(n2720));
sg13g2_nor2_2 U2792 (.A(n4165), .B(n653), .Y(n2722));
sg13g2_inv_4 U2793 (.A(n2721), .Y(n2715));
sg13g2_o21ai_1 U2794 (.A1(n4325), .A2(n2719), .B1(n2723), .Y(n2721));
sg13g2_a21oi_2 U2795 (.A1(data_i_57_), .A2(n4308), .B1(n2724), .Y(n2723));
sg13g2_nor2_2 U2796 (.A(n555), .B(n653), .Y(n2724));
sg13g2_inv_4 U2797 (.A(mixcol_data_o_57), .Y(n653));
sg13g2_inv_4 U2798 (.A(subbytes_data_o_57), .Y(n2719));
sg13g2_a21oi_2 U2800 (.A1(n4313), .A2(n2727), .B1(n2728), .Y(n2726));
sg13g2_nor2_2 U2801 (.A(n2729), .B(n4310), .Y(n2728));
sg13g2_o21ai_1 U2802 (.A1(n4167), .A2(n2729), .B1(n2730), .Y(n2727));
sg13g2_a21oi_2 U2803 (.A1(n4315), .A2(n2731), .B1(n2732), .Y(n2730));
sg13g2_nor2_2 U2804 (.A(n4164), .B(n655), .Y(n2732));
sg13g2_inv_4 U2805 (.A(n2731), .Y(n2725));
sg13g2_o21ai_1 U2806 (.A1(n4330), .A2(n2729), .B1(n2733), .Y(n2731));
sg13g2_a21oi_2 U2807 (.A1(data_i_56_), .A2(n4308), .B1(n2734), .Y(n2733));
sg13g2_nor2_2 U2808 (.A(n555), .B(n655), .Y(n2734));
sg13g2_inv_4 U2809 (.A(mixcol_data_o_56), .Y(n655));
sg13g2_inv_4 U2810 (.A(subbytes_data_o_56), .Y(n2729));
sg13g2_a21oi_2 U2812 (.A1(n4312), .A2(n2737), .B1(n2738), .Y(n2736));
sg13g2_nor2_2 U2813 (.A(n2739), .B(n2248), .Y(n2738));
sg13g2_o21ai_1 U2814 (.A1(n553), .A2(n2739), .B1(n2740), .Y(n2737));
sg13g2_a21oi_2 U2815 (.A1(n4315), .A2(n2741), .B1(n2742), .Y(n2740));
sg13g2_nor2_2 U2816 (.A(n4165), .B(n657), .Y(n2742));
sg13g2_inv_4 U2817 (.A(n2741), .Y(n2735));
sg13g2_o21ai_1 U2818 (.A1(n4329), .A2(n2739), .B1(n2743), .Y(n2741));
sg13g2_a21oi_2 U2819 (.A1(data_i_55_), .A2(n4308), .B1(n2744), .Y(n2743));
sg13g2_nor2_2 U2820 (.A(n555), .B(n657), .Y(n2744));
sg13g2_inv_4 U2821 (.A(mixcol_data_o_55), .Y(n657));
sg13g2_inv_4 U2822 (.A(subbytes_data_o_55), .Y(n2739));
sg13g2_a21oi_2 U2824 (.A1(n4313), .A2(n2747), .B1(n2748), .Y(n2746));
sg13g2_nor2_2 U2825 (.A(n2749), .B(n4310), .Y(n2748));
sg13g2_o21ai_1 U2826 (.A1(n4167), .A2(n2749), .B1(n2750), .Y(n2747));
sg13g2_a21oi_2 U2827 (.A1(n4315), .A2(n2751), .B1(n2752), .Y(n2750));
sg13g2_nor2_2 U2828 (.A(n4164), .B(n659), .Y(n2752));
sg13g2_inv_4 U2829 (.A(n2751), .Y(n2745));
sg13g2_o21ai_1 U2830 (.A1(n4330), .A2(n2749), .B1(n2753), .Y(n2751));
sg13g2_a21oi_2 U2831 (.A1(data_i_54_), .A2(n4308), .B1(n2754), .Y(n2753));
sg13g2_nor2_2 U2832 (.A(n555), .B(n659), .Y(n2754));
sg13g2_inv_4 U2833 (.A(mixcol_data_o_54), .Y(n659));
sg13g2_inv_4 U2834 (.A(subbytes_data_o_54), .Y(n2749));
sg13g2_a21oi_2 U2836 (.A1(n4312), .A2(n2757), .B1(n2758), .Y(n2756));
sg13g2_nor2_2 U2837 (.A(n2759), .B(n4310), .Y(n2758));
sg13g2_o21ai_1 U2838 (.A1(n553), .A2(n2759), .B1(n2760), .Y(n2757));
sg13g2_a21oi_2 U2839 (.A1(n4315), .A2(n2761), .B1(n2762), .Y(n2760));
sg13g2_nor2_2 U2840 (.A(n4164), .B(n661), .Y(n2762));
sg13g2_inv_4 U2841 (.A(n2761), .Y(n2755));
sg13g2_o21ai_1 U2842 (.A1(n4326), .A2(n2759), .B1(n2763), .Y(n2761));
sg13g2_a21oi_2 U2843 (.A1(data_i_53_), .A2(n4307), .B1(n2764), .Y(n2763));
sg13g2_nor2_2 U2844 (.A(n555), .B(n661), .Y(n2764));
sg13g2_inv_4 U2845 (.A(mixcol_data_o_53), .Y(n661));
sg13g2_inv_4 U2846 (.A(subbytes_data_o_53), .Y(n2759));
sg13g2_a21oi_2 U2848 (.A1(n4313), .A2(n2767), .B1(n2768), .Y(n2766));
sg13g2_nor2_2 U2849 (.A(n2769), .B(n4310), .Y(n2768));
sg13g2_o21ai_1 U2850 (.A1(n553), .A2(n2769), .B1(n2770), .Y(n2767));
sg13g2_a21oi_2 U2851 (.A1(n4315), .A2(n2771), .B1(n2772), .Y(n2770));
sg13g2_nor2_2 U2852 (.A(n4164), .B(n663), .Y(n2772));
sg13g2_inv_4 U2853 (.A(n2771), .Y(n2765));
sg13g2_o21ai_1 U2854 (.A1(n4330), .A2(n2769), .B1(n2773), .Y(n2771));
sg13g2_a21oi_2 U2855 (.A1(data_i_52_), .A2(n4307), .B1(n2774), .Y(n2773));
sg13g2_nor2_2 U2856 (.A(n555), .B(n663), .Y(n2774));
sg13g2_inv_4 U2857 (.A(mixcol_data_o_52), .Y(n663));
sg13g2_inv_4 U2858 (.A(subbytes_data_o_52), .Y(n2769));
sg13g2_a21oi_2 U2860 (.A1(n4312), .A2(n2777), .B1(n2778), .Y(n2776));
sg13g2_nor2_2 U2861 (.A(n2779), .B(n4310), .Y(n2778));
sg13g2_o21ai_1 U2862 (.A1(n4167), .A2(n2779), .B1(n2780), .Y(n2777));
sg13g2_a21oi_2 U2863 (.A1(n4315), .A2(n2781), .B1(n2782), .Y(n2780));
sg13g2_nor2_2 U2864 (.A(n4165), .B(n665), .Y(n2782));
sg13g2_inv_4 U2865 (.A(n2781), .Y(n2775));
sg13g2_o21ai_1 U2866 (.A1(n4327), .A2(n2779), .B1(n2783), .Y(n2781));
sg13g2_a21oi_2 U2867 (.A1(data_i_51_), .A2(n4308), .B1(n2784), .Y(n2783));
sg13g2_nor2_2 U2868 (.A(n555), .B(n665), .Y(n2784));
sg13g2_inv_4 U2869 (.A(mixcol_data_o_51), .Y(n665));
sg13g2_inv_4 U2870 (.A(subbytes_data_o_51), .Y(n2779));
sg13g2_a21oi_2 U2872 (.A1(n4312), .A2(n2787), .B1(n2788), .Y(n2786));
sg13g2_nor2_2 U2873 (.A(n2789), .B(n4310), .Y(n2788));
sg13g2_o21ai_1 U2874 (.A1(n4167), .A2(n2789), .B1(n2790), .Y(n2787));
sg13g2_a21oi_2 U2875 (.A1(n4315), .A2(n2791), .B1(n2792), .Y(n2790));
sg13g2_nor2_2 U2876 (.A(n4165), .B(n667), .Y(n2792));
sg13g2_inv_4 U2877 (.A(n2791), .Y(n2785));
sg13g2_o21ai_1 U2878 (.A1(n4326), .A2(n2789), .B1(n2793), .Y(n2791));
sg13g2_a21oi_2 U2879 (.A1(data_i_50_), .A2(n4308), .B1(n2794), .Y(n2793));
sg13g2_nor2_2 U2880 (.A(n555), .B(n667), .Y(n2794));
sg13g2_inv_4 U2881 (.A(mixcol_data_o_50), .Y(n667));
sg13g2_inv_4 U2882 (.A(subbytes_data_o_50), .Y(n2789));
sg13g2_a21oi_2 U2884 (.A1(n4312), .A2(n2797), .B1(n2798), .Y(n2796));
sg13g2_nor2_2 U2885 (.A(n2799), .B(n4310), .Y(n2798));
sg13g2_o21ai_1 U2886 (.A1(n553), .A2(n2799), .B1(n2800), .Y(n2797));
sg13g2_a21oi_2 U2887 (.A1(n4315), .A2(n2801), .B1(n2802), .Y(n2800));
sg13g2_nor2_2 U2888 (.A(n4164), .B(n669), .Y(n2802));
sg13g2_inv_4 U2889 (.A(n2801), .Y(n2795));
sg13g2_o21ai_1 U2890 (.A1(n4329), .A2(n2799), .B1(n2803), .Y(n2801));
sg13g2_a21oi_2 U2891 (.A1(data_i_4_), .A2(n4307), .B1(n2804), .Y(n2803));
sg13g2_nor2_2 U2892 (.A(n555), .B(n669), .Y(n2804));
sg13g2_inv_4 U2893 (.A(mixcol_data_o_4), .Y(n669));
sg13g2_inv_4 U2894 (.A(subbytes_data_o_4), .Y(n2799));
sg13g2_a21oi_2 U2896 (.A1(n4312), .A2(n2807), .B1(n2808), .Y(n2806));
sg13g2_nor2_2 U2897 (.A(n2809), .B(n4310), .Y(n2808));
sg13g2_o21ai_1 U2898 (.A1(n4167), .A2(n2809), .B1(n2810), .Y(n2807));
sg13g2_a21oi_2 U2899 (.A1(n4315), .A2(n2811), .B1(n2812), .Y(n2810));
sg13g2_nor2_2 U2900 (.A(n4164), .B(n671), .Y(n2812));
sg13g2_inv_4 U2901 (.A(n2811), .Y(n2805));
sg13g2_o21ai_1 U2902 (.A1(n4330), .A2(n2809), .B1(n2813), .Y(n2811));
sg13g2_a21oi_2 U2903 (.A1(data_i_49_), .A2(n4308), .B1(n2814), .Y(n2813));
sg13g2_nor2_2 U2904 (.A(n555), .B(n671), .Y(n2814));
sg13g2_inv_4 U2905 (.A(mixcol_data_o_49), .Y(n671));
sg13g2_inv_4 U2906 (.A(subbytes_data_o_49), .Y(n2809));
sg13g2_a21oi_2 U2908 (.A1(n4313), .A2(n2817), .B1(n2818), .Y(n2816));
sg13g2_nor2_2 U2909 (.A(n2819), .B(n4310), .Y(n2818));
sg13g2_o21ai_1 U2910 (.A1(n553), .A2(n2819), .B1(n2820), .Y(n2817));
sg13g2_a21oi_2 U2911 (.A1(n4315), .A2(n2821), .B1(n2822), .Y(n2820));
sg13g2_nor2_2 U2912 (.A(n4165), .B(n673), .Y(n2822));
sg13g2_inv_4 U2913 (.A(n2821), .Y(n2815));
sg13g2_o21ai_1 U2914 (.A1(n4327), .A2(n2819), .B1(n2823), .Y(n2821));
sg13g2_a21oi_2 U2915 (.A1(data_i_48_), .A2(n4307), .B1(n2824), .Y(n2823));
sg13g2_nor2_2 U2916 (.A(n555), .B(n673), .Y(n2824));
sg13g2_inv_4 U2917 (.A(mixcol_data_o_48), .Y(n673));
sg13g2_inv_4 U2918 (.A(subbytes_data_o_48), .Y(n2819));
sg13g2_o21ai_1 U2919 (.A1(state), .A2(n2825), .B1(n2826), .Y(addroundkey_data_i_47));
sg13g2_a21oi_2 U2920 (.A1(n2244), .A2(n2827), .B1(n2828), .Y(n2826));
sg13g2_nor2_2 U2921 (.A(n2829), .B(n4310), .Y(n2828));
sg13g2_o21ai_1 U2922 (.A1(n4167), .A2(n2829), .B1(n2830), .Y(n2827));
sg13g2_a21oi_2 U2923 (.A1(n4315), .A2(n2831), .B1(n2832), .Y(n2830));
sg13g2_nor2_2 U2924 (.A(n4164), .B(n675), .Y(n2832));
sg13g2_inv_4 U2925 (.A(n2831), .Y(n2825));
sg13g2_o21ai_1 U2926 (.A1(n4330), .A2(n2829), .B1(n2833), .Y(n2831));
sg13g2_a21oi_2 U2927 (.A1(data_i_47_), .A2(n4307), .B1(n2834), .Y(n2833));
sg13g2_nor2_2 U2928 (.A(n555), .B(n675), .Y(n2834));
sg13g2_inv_4 U2929 (.A(mixcol_data_o_47), .Y(n675));
sg13g2_inv_4 U2930 (.A(subbytes_data_o_47), .Y(n2829));
sg13g2_a21oi_2 U2932 (.A1(n2244), .A2(n2837), .B1(n2838), .Y(n2836));
sg13g2_nor2_2 U2933 (.A(n2839), .B(n4310), .Y(n2838));
sg13g2_o21ai_1 U2934 (.A1(n553), .A2(n2839), .B1(n2840), .Y(n2837));
sg13g2_a21oi_2 U2935 (.A1(n4315), .A2(n2841), .B1(n2842), .Y(n2840));
sg13g2_nor2_2 U2936 (.A(n4164), .B(n677), .Y(n2842));
sg13g2_inv_4 U2937 (.A(n2841), .Y(n2835));
sg13g2_o21ai_1 U2938 (.A1(n4328), .A2(n2839), .B1(n2843), .Y(n2841));
sg13g2_a21oi_2 U2939 (.A1(data_i_46_), .A2(n4307), .B1(n2844), .Y(n2843));
sg13g2_nor2_2 U2940 (.A(n555), .B(n677), .Y(n2844));
sg13g2_inv_4 U2941 (.A(mixcol_data_o_46), .Y(n677));
sg13g2_inv_4 U2942 (.A(subbytes_data_o_46), .Y(n2839));
sg13g2_a21oi_2 U2944 (.A1(n4313), .A2(n2847), .B1(n2848), .Y(n2846));
sg13g2_nor2_2 U2945 (.A(n2849), .B(n4310), .Y(n2848));
sg13g2_o21ai_1 U2946 (.A1(n4167), .A2(n2849), .B1(n2850), .Y(n2847));
sg13g2_a21oi_2 U2947 (.A1(n4315), .A2(n2851), .B1(n2852), .Y(n2850));
sg13g2_nor2_2 U2948 (.A(n4164), .B(n679), .Y(n2852));
sg13g2_inv_4 U2949 (.A(n2851), .Y(n2845));
sg13g2_o21ai_1 U2950 (.A1(n4328), .A2(n2849), .B1(n2853), .Y(n2851));
sg13g2_a21oi_2 U2951 (.A1(data_i_45_), .A2(n4307), .B1(n2854), .Y(n2853));
sg13g2_nor2_2 U2952 (.A(n555), .B(n679), .Y(n2854));
sg13g2_inv_4 U2953 (.A(mixcol_data_o_45), .Y(n679));
sg13g2_inv_4 U2954 (.A(subbytes_data_o_45), .Y(n2849));
sg13g2_a21oi_2 U2956 (.A1(n4313), .A2(n2857), .B1(n2858), .Y(n2856));
sg13g2_nor2_2 U2957 (.A(n2859), .B(n4310), .Y(n2858));
sg13g2_o21ai_1 U2958 (.A1(n4167), .A2(n2859), .B1(n2860), .Y(n2857));
sg13g2_a21oi_2 U2959 (.A1(n4315), .A2(n2861), .B1(n2862), .Y(n2860));
sg13g2_nor2_2 U2960 (.A(n4165), .B(n681), .Y(n2862));
sg13g2_inv_4 U2961 (.A(n2861), .Y(n2855));
sg13g2_o21ai_1 U2962 (.A1(n4330), .A2(n2859), .B1(n2863), .Y(n2861));
sg13g2_a21oi_2 U2963 (.A1(data_i_44_), .A2(n4307), .B1(n2864), .Y(n2863));
sg13g2_nor2_2 U2964 (.A(n555), .B(n681), .Y(n2864));
sg13g2_inv_4 U2965 (.A(mixcol_data_o_44), .Y(n681));
sg13g2_inv_4 U2966 (.A(subbytes_data_o_44), .Y(n2859));
sg13g2_a21oi_2 U2968 (.A1(n2244), .A2(n2867), .B1(n2868), .Y(n2866));
sg13g2_nor2_2 U2969 (.A(n2869), .B(n2248), .Y(n2868));
sg13g2_o21ai_1 U2970 (.A1(n553), .A2(n2869), .B1(n2870), .Y(n2867));
sg13g2_a21oi_2 U2971 (.A1(n4315), .A2(n2871), .B1(n2872), .Y(n2870));
sg13g2_nor2_2 U2972 (.A(n4164), .B(n683), .Y(n2872));
sg13g2_inv_4 U2973 (.A(n2871), .Y(n2865));
sg13g2_o21ai_1 U2974 (.A1(n4326), .A2(n2869), .B1(n2873), .Y(n2871));
sg13g2_a21oi_2 U2975 (.A1(data_i_43_), .A2(n4307), .B1(n2874), .Y(n2873));
sg13g2_nor2_2 U2976 (.A(n555), .B(n683), .Y(n2874));
sg13g2_inv_4 U2977 (.A(mixcol_data_o_43), .Y(n683));
sg13g2_inv_4 U2978 (.A(subbytes_data_o_43), .Y(n2869));
sg13g2_a21oi_2 U2980 (.A1(n4313), .A2(n2877), .B1(n2878), .Y(n2876));
sg13g2_nor2_2 U2981 (.A(n2879), .B(n2248), .Y(n2878));
sg13g2_o21ai_1 U2982 (.A1(n553), .A2(n2879), .B1(n2880), .Y(n2877));
sg13g2_a21oi_2 U2983 (.A1(n4315), .A2(n2881), .B1(n2882), .Y(n2880));
sg13g2_nor2_2 U2984 (.A(n4165), .B(n685), .Y(n2882));
sg13g2_inv_4 U2985 (.A(n2881), .Y(n2875));
sg13g2_o21ai_1 U2986 (.A1(n4327), .A2(n2879), .B1(n2883), .Y(n2881));
sg13g2_a21oi_2 U2987 (.A1(data_i_42_), .A2(n4307), .B1(n2884), .Y(n2883));
sg13g2_nor2_2 U2988 (.A(n555), .B(n685), .Y(n2884));
sg13g2_inv_4 U2989 (.A(mixcol_data_o_42), .Y(n685));
sg13g2_inv_4 U2990 (.A(subbytes_data_o_42), .Y(n2879));
sg13g2_a21oi_2 U2992 (.A1(n2244), .A2(n2887), .B1(n2888), .Y(n2886));
sg13g2_nor2_2 U2993 (.A(n2889), .B(n2248), .Y(n2888));
sg13g2_o21ai_1 U2994 (.A1(n553), .A2(n2889), .B1(n2890), .Y(n2887));
sg13g2_a21oi_2 U2995 (.A1(n4315), .A2(n2891), .B1(n2892), .Y(n2890));
sg13g2_nor2_2 U2996 (.A(n4164), .B(n687), .Y(n2892));
sg13g2_inv_4 U2997 (.A(n2891), .Y(n2885));
sg13g2_o21ai_1 U2998 (.A1(n4330), .A2(n2889), .B1(n2893), .Y(n2891));
sg13g2_a21oi_2 U2999 (.A1(data_i_41_), .A2(n4307), .B1(n2894), .Y(n2893));
sg13g2_nor2_2 U3000 (.A(n555), .B(n687), .Y(n2894));
sg13g2_inv_4 U3001 (.A(mixcol_data_o_41), .Y(n687));
sg13g2_inv_4 U3002 (.A(subbytes_data_o_41), .Y(n2889));
sg13g2_a21oi_2 U3004 (.A1(n4313), .A2(n2897), .B1(n2898), .Y(n2896));
sg13g2_nor2_2 U3005 (.A(n2899), .B(n2248), .Y(n2898));
sg13g2_o21ai_1 U3006 (.A1(n4167), .A2(n2899), .B1(n2900), .Y(n2897));
sg13g2_a21oi_2 U3007 (.A1(n4315), .A2(n2901), .B1(n2902), .Y(n2900));
sg13g2_nor2_2 U3008 (.A(n4165), .B(n689), .Y(n2902));
sg13g2_inv_4 U3009 (.A(n2901), .Y(n2895));
sg13g2_o21ai_1 U3010 (.A1(n4329), .A2(n2899), .B1(n2903), .Y(n2901));
sg13g2_a21oi_2 U3011 (.A1(data_i_40_), .A2(n4307), .B1(n2904), .Y(n2903));
sg13g2_nor2_2 U3012 (.A(n555), .B(n689), .Y(n2904));
sg13g2_inv_4 U3013 (.A(mixcol_data_o_40), .Y(n689));
sg13g2_inv_4 U3014 (.A(subbytes_data_o_40), .Y(n2899));
sg13g2_a21oi_2 U3016 (.A1(n4312), .A2(n2907), .B1(n2908), .Y(n2906));
sg13g2_nor2_2 U3017 (.A(n2909), .B(n2248), .Y(n2908));
sg13g2_o21ai_1 U3018 (.A1(n4167), .A2(n2909), .B1(n2910), .Y(n2907));
sg13g2_a21oi_2 U3019 (.A1(n4315), .A2(n2911), .B1(n2912), .Y(n2910));
sg13g2_nor2_2 U3020 (.A(n4165), .B(n691), .Y(n2912));
sg13g2_inv_4 U3021 (.A(n2911), .Y(n2905));
sg13g2_o21ai_1 U3022 (.A1(n4328), .A2(n2909), .B1(n2913), .Y(n2911));
sg13g2_a21oi_2 U3023 (.A1(data_i_3_), .A2(n4307), .B1(n2914), .Y(n2913));
sg13g2_nor2_2 U3024 (.A(n555), .B(n691), .Y(n2914));
sg13g2_inv_4 U3025 (.A(mixcol_data_o_3), .Y(n691));
sg13g2_inv_4 U3026 (.A(subbytes_data_o_3), .Y(n2909));
sg13g2_nor2_2 U3029 (.A(n2919), .B(n2248), .Y(n2918));
sg13g2_o21ai_1 U3030 (.A1(n4167), .A2(n2919), .B1(n2920), .Y(n2917));
sg13g2_a21oi_2 U3031 (.A1(n4315), .A2(n2921), .B1(n2922), .Y(n2920));
sg13g2_nor2_2 U3032 (.A(n4164), .B(n693), .Y(n2922));
sg13g2_inv_4 U3033 (.A(n2921), .Y(n2915));
sg13g2_o21ai_1 U3034 (.A1(n4326), .A2(n2919), .B1(n2923), .Y(n2921));
sg13g2_a21oi_2 U3035 (.A1(data_i_39_), .A2(n4307), .B1(n2924), .Y(n2923));
sg13g2_nor2_2 U3036 (.A(n555), .B(n693), .Y(n2924));
sg13g2_inv_4 U3037 (.A(mixcol_data_o_39), .Y(n693));
sg13g2_inv_4 U3038 (.A(subbytes_data_o_39), .Y(n2919));
sg13g2_a21oi_2 U3040 (.A1(n4313), .A2(n2927), .B1(n2928), .Y(n2926));
sg13g2_nor2_2 U3041 (.A(n2929), .B(n2248), .Y(n2928));
sg13g2_o21ai_1 U3042 (.A1(n553), .A2(n2929), .B1(n2930), .Y(n2927));
sg13g2_a21oi_2 U3043 (.A1(n4315), .A2(n2931), .B1(n2932), .Y(n2930));
sg13g2_nor2_2 U3044 (.A(n4164), .B(n695), .Y(n2932));
sg13g2_inv_4 U3045 (.A(n2931), .Y(n2925));
sg13g2_o21ai_1 U3046 (.A1(n4325), .A2(n2929), .B1(n2933), .Y(n2931));
sg13g2_nor2_2 U3048 (.A(n555), .B(n695), .Y(n2934));
sg13g2_inv_4 U3049 (.A(mixcol_data_o_38), .Y(n695));
sg13g2_inv_4 U3050 (.A(subbytes_data_o_38), .Y(n2929));
sg13g2_a21oi_2 U3052 (.A1(n4313), .A2(n2937), .B1(n2938), .Y(n2936));
sg13g2_nor2_2 U3053 (.A(n2939), .B(n2248), .Y(n2938));
sg13g2_o21ai_1 U3054 (.A1(n553), .A2(n2939), .B1(n2940), .Y(n2937));
sg13g2_a21oi_2 U3055 (.A1(n4315), .A2(n2941), .B1(n2942), .Y(n2940));
sg13g2_nor2_2 U3056 (.A(n4165), .B(n697), .Y(n2942));
sg13g2_inv_4 U3057 (.A(n2941), .Y(n2935));
sg13g2_o21ai_1 U3058 (.A1(n4330), .A2(n2939), .B1(n2943), .Y(n2941));
sg13g2_nor2_2 U3060 (.A(n555), .B(n697), .Y(n2944));
sg13g2_inv_4 U3061 (.A(mixcol_data_o_37), .Y(n697));
sg13g2_inv_4 U3062 (.A(subbytes_data_o_37), .Y(n2939));
sg13g2_a21oi_2 U3064 (.A1(n4313), .A2(n2947), .B1(n2948), .Y(n2946));
sg13g2_nor2_2 U3065 (.A(n2949), .B(n2248), .Y(n2948));
sg13g2_o21ai_1 U3066 (.A1(n553), .A2(n2949), .B1(n2950), .Y(n2947));
sg13g2_a21oi_2 U3067 (.A1(n4315), .A2(n2951), .B1(n2952), .Y(n2950));
sg13g2_nor2_2 U3068 (.A(n4164), .B(n699), .Y(n2952));
sg13g2_inv_4 U3069 (.A(n2951), .Y(n2945));
sg13g2_o21ai_1 U3070 (.A1(n4330), .A2(n2949), .B1(n2953), .Y(n2951));
sg13g2_a21oi_2 U3071 (.A1(data_i_36_), .A2(n4308), .B1(n2954), .Y(n2953));
sg13g2_nor2_2 U3072 (.A(n555), .B(n699), .Y(n2954));
sg13g2_inv_4 U3073 (.A(mixcol_data_o_36), .Y(n699));
sg13g2_inv_4 U3074 (.A(subbytes_data_o_36), .Y(n2949));
sg13g2_a21oi_2 U3076 (.A1(n4313), .A2(n2957), .B1(n2958), .Y(n2956));
sg13g2_nor2_2 U3077 (.A(n2959), .B(n2248), .Y(n2958));
sg13g2_o21ai_1 U3078 (.A1(n4167), .A2(n2959), .B1(n2960), .Y(n2957));
sg13g2_a21oi_2 U3079 (.A1(n4315), .A2(n2961), .B1(n2962), .Y(n2960));
sg13g2_nor2_2 U3080 (.A(n4165), .B(n701), .Y(n2962));
sg13g2_inv_4 U3081 (.A(n2961), .Y(n2955));
sg13g2_o21ai_1 U3082 (.A1(n4325), .A2(n2959), .B1(n2963), .Y(n2961));
sg13g2_a21oi_2 U3083 (.A1(data_i_35_), .A2(n4307), .B1(n2964), .Y(n2963));
sg13g2_nor2_2 U3084 (.A(n555), .B(n701), .Y(n2964));
sg13g2_inv_4 U3085 (.A(mixcol_data_o_35), .Y(n701));
sg13g2_inv_4 U3086 (.A(subbytes_data_o_35), .Y(n2959));
sg13g2_a21oi_2 U3088 (.A1(n4313), .A2(n2967), .B1(n2968), .Y(n2966));
sg13g2_nor2_2 U3089 (.A(n2969), .B(n2248), .Y(n2968));
sg13g2_o21ai_1 U3090 (.A1(n4167), .A2(n2969), .B1(n2970), .Y(n2967));
sg13g2_a21oi_2 U3091 (.A1(n4315), .A2(n2971), .B1(n2972), .Y(n2970));
sg13g2_nor2_2 U3092 (.A(n4164), .B(n703), .Y(n2972));
sg13g2_inv_4 U3093 (.A(n2971), .Y(n2965));
sg13g2_o21ai_1 U3094 (.A1(n4330), .A2(n2969), .B1(n2973), .Y(n2971));
sg13g2_a21oi_2 U3095 (.A1(data_i_34_), .A2(n4308), .B1(n2974), .Y(n2973));
sg13g2_nor2_2 U3096 (.A(n555), .B(n703), .Y(n2974));
sg13g2_inv_4 U3097 (.A(mixcol_data_o_34), .Y(n703));
sg13g2_inv_4 U3098 (.A(subbytes_data_o_34), .Y(n2969));
sg13g2_a21oi_2 U3100 (.A1(n4313), .A2(n2977), .B1(n2978), .Y(n2976));
sg13g2_nor2_2 U3101 (.A(n2979), .B(n2248), .Y(n2978));
sg13g2_o21ai_1 U3102 (.A1(n4167), .A2(n2979), .B1(n2980), .Y(n2977));
sg13g2_a21oi_2 U3103 (.A1(n4315), .A2(n2981), .B1(n2982), .Y(n2980));
sg13g2_nor2_2 U3104 (.A(n4165), .B(n705), .Y(n2982));
sg13g2_inv_4 U3105 (.A(n2981), .Y(n2975));
sg13g2_o21ai_1 U3106 (.A1(n4329), .A2(n2979), .B1(n2983), .Y(n2981));
sg13g2_a21oi_2 U3107 (.A1(data_i_33_), .A2(n4307), .B1(n2984), .Y(n2983));
sg13g2_nor2_2 U3108 (.A(n555), .B(n705), .Y(n2984));
sg13g2_inv_4 U3109 (.A(mixcol_data_o_33), .Y(n705));
sg13g2_inv_4 U3110 (.A(subbytes_data_o_33), .Y(n2979));
sg13g2_a21oi_2 U3112 (.A1(n4313), .A2(n2987), .B1(n2988), .Y(n2986));
sg13g2_nor2_2 U3113 (.A(n2989), .B(n4310), .Y(n2988));
sg13g2_o21ai_1 U3114 (.A1(n4167), .A2(n2989), .B1(n2990), .Y(n2987));
sg13g2_a21oi_2 U3115 (.A1(n4315), .A2(n2991), .B1(n2992), .Y(n2990));
sg13g2_nor2_2 U3116 (.A(n4164), .B(n707), .Y(n2992));
sg13g2_inv_4 U3117 (.A(n2991), .Y(n2985));
sg13g2_o21ai_1 U3118 (.A1(n4330), .A2(n2989), .B1(n2993), .Y(n2991));
sg13g2_a21oi_2 U3119 (.A1(data_i_32_), .A2(n4308), .B1(n2994), .Y(n2993));
sg13g2_nor2_2 U3120 (.A(n555), .B(n707), .Y(n2994));
sg13g2_inv_4 U3121 (.A(mixcol_data_o_32), .Y(n707));
sg13g2_inv_4 U3122 (.A(subbytes_data_o_32), .Y(n2989));
sg13g2_a21oi_2 U3124 (.A1(n4313), .A2(n2997), .B1(n2998), .Y(n2996));
sg13g2_nor2_2 U3125 (.A(n2999), .B(n2248), .Y(n2998));
sg13g2_o21ai_1 U3126 (.A1(n553), .A2(n2999), .B1(n3000), .Y(n2997));
sg13g2_a21oi_2 U3127 (.A1(n4315), .A2(n3001), .B1(n3002), .Y(n3000));
sg13g2_nor2_2 U3128 (.A(n4165), .B(n709), .Y(n3002));
sg13g2_inv_4 U3129 (.A(n3001), .Y(n2995));
sg13g2_o21ai_1 U3130 (.A1(n4328), .A2(n2999), .B1(n3003), .Y(n3001));
sg13g2_a21oi_2 U3131 (.A1(data_i_31_), .A2(n4308), .B1(n3004), .Y(n3003));
sg13g2_nor2_2 U3132 (.A(n555), .B(n709), .Y(n3004));
sg13g2_inv_4 U3133 (.A(mixcol_data_o_31), .Y(n709));
sg13g2_inv_4 U3134 (.A(subbytes_data_o_31), .Y(n2999));
sg13g2_a21oi_2 U3136 (.A1(n4313), .A2(n3007), .B1(n3008), .Y(n3006));
sg13g2_nor2_2 U3137 (.A(n3009), .B(n4310), .Y(n3008));
sg13g2_o21ai_1 U3138 (.A1(n553), .A2(n3009), .B1(n3010), .Y(n3007));
sg13g2_a21oi_2 U3139 (.A1(n4315), .A2(n3011), .B1(n3012), .Y(n3010));
sg13g2_nor2_2 U3140 (.A(n4164), .B(n711), .Y(n3012));
sg13g2_inv_4 U3141 (.A(n3011), .Y(n3005));
sg13g2_o21ai_1 U3142 (.A1(n4325), .A2(n3009), .B1(n3013), .Y(n3011));
sg13g2_a21oi_2 U3143 (.A1(data_i_30_), .A2(n4308), .B1(n3014), .Y(n3013));
sg13g2_nor2_2 U3144 (.A(n555), .B(n711), .Y(n3014));
sg13g2_inv_4 U3145 (.A(mixcol_data_o_30), .Y(n711));
sg13g2_inv_4 U3146 (.A(subbytes_data_o_30), .Y(n3009));
sg13g2_a21oi_2 U3148 (.A1(n4313), .A2(n3017), .B1(n3018), .Y(n3016));
sg13g2_nor2_2 U3149 (.A(n3019), .B(n2248), .Y(n3018));
sg13g2_o21ai_1 U3150 (.A1(n553), .A2(n3019), .B1(n3020), .Y(n3017));
sg13g2_a21oi_2 U3151 (.A1(n4315), .A2(n3021), .B1(n3022), .Y(n3020));
sg13g2_nor2_2 U3152 (.A(n4164), .B(n713), .Y(n3022));
sg13g2_inv_4 U3153 (.A(n3021), .Y(n3015));
sg13g2_o21ai_1 U3154 (.A1(n4330), .A2(n3019), .B1(n3023), .Y(n3021));
sg13g2_a21oi_2 U3155 (.A1(data_i_2_), .A2(n4308), .B1(n3024), .Y(n3023));
sg13g2_nor2_2 U3156 (.A(n555), .B(n713), .Y(n3024));
sg13g2_inv_4 U3157 (.A(mixcol_data_o_2), .Y(n713));
sg13g2_inv_4 U3158 (.A(subbytes_data_o_2), .Y(n3019));
sg13g2_a21oi_2 U3160 (.A1(n4313), .A2(n3027), .B1(n3028), .Y(n3026));
sg13g2_nor2_2 U3161 (.A(n3029), .B(n2248), .Y(n3028));
sg13g2_o21ai_1 U3162 (.A1(n553), .A2(n3029), .B1(n3030), .Y(n3027));
sg13g2_a21oi_2 U3163 (.A1(n4315), .A2(n3031), .B1(n3032), .Y(n3030));
sg13g2_nor2_2 U3164 (.A(n4164), .B(n715), .Y(n3032));
sg13g2_inv_4 U3165 (.A(n3031), .Y(n3025));
sg13g2_o21ai_1 U3166 (.A1(n4327), .A2(n3029), .B1(n3033), .Y(n3031));
sg13g2_a21oi_2 U3167 (.A1(data_i_29_), .A2(n4307), .B1(n3034), .Y(n3033));
sg13g2_nor2_2 U3168 (.A(n555), .B(n715), .Y(n3034));
sg13g2_inv_4 U3169 (.A(mixcol_data_o_29), .Y(n715));
sg13g2_inv_4 U3170 (.A(subbytes_data_o_29), .Y(n3029));
sg13g2_a21oi_2 U3172 (.A1(n4312), .A2(n3037), .B1(n3038), .Y(n3036));
sg13g2_nor2_2 U3173 (.A(n3039), .B(n2248), .Y(n3038));
sg13g2_o21ai_1 U3174 (.A1(n4167), .A2(n3039), .B1(n3040), .Y(n3037));
sg13g2_a21oi_2 U3175 (.A1(n4315), .A2(n3041), .B1(n3042), .Y(n3040));
sg13g2_nor2_2 U3176 (.A(n4164), .B(n717), .Y(n3042));
sg13g2_inv_4 U3177 (.A(n3041), .Y(n3035));
sg13g2_o21ai_1 U3178 (.A1(n4329), .A2(n3039), .B1(n3043), .Y(n3041));
sg13g2_a21oi_2 U3179 (.A1(data_i_28_), .A2(n4307), .B1(n3044), .Y(n3043));
sg13g2_nor2_2 U3180 (.A(n555), .B(n717), .Y(n3044));
sg13g2_inv_4 U3181 (.A(mixcol_data_o_28), .Y(n717));
sg13g2_inv_4 U3182 (.A(subbytes_data_o_28), .Y(n3039));
sg13g2_a21oi_2 U3184 (.A1(n4312), .A2(n3047), .B1(n3048), .Y(n3046));
sg13g2_nor2_2 U3185 (.A(n3049), .B(n2248), .Y(n3048));
sg13g2_o21ai_1 U3186 (.A1(n4167), .A2(n3049), .B1(n3050), .Y(n3047));
sg13g2_a21oi_2 U3187 (.A1(n4315), .A2(n3051), .B1(n3052), .Y(n3050));
sg13g2_nor2_2 U3188 (.A(n4165), .B(n719), .Y(n3052));
sg13g2_inv_4 U3189 (.A(n3051), .Y(n3045));
sg13g2_o21ai_1 U3190 (.A1(n4330), .A2(n3049), .B1(n3053), .Y(n3051));
sg13g2_a21oi_2 U3191 (.A1(data_i_27_), .A2(n4307), .B1(n3054), .Y(n3053));
sg13g2_nor2_2 U3192 (.A(n555), .B(n719), .Y(n3054));
sg13g2_inv_4 U3193 (.A(mixcol_data_o_27), .Y(n719));
sg13g2_inv_4 U3194 (.A(subbytes_data_o_27), .Y(n3049));
sg13g2_a21oi_2 U3196 (.A1(n4313), .A2(n3057), .B1(n3058), .Y(n3056));
sg13g2_nor2_2 U3197 (.A(n3059), .B(n2248), .Y(n3058));
sg13g2_o21ai_1 U3198 (.A1(n4167), .A2(n3059), .B1(n3060), .Y(n3057));
sg13g2_a21oi_2 U3199 (.A1(n4315), .A2(n3061), .B1(n3062), .Y(n3060));
sg13g2_nor2_2 U3200 (.A(n4165), .B(n721), .Y(n3062));
sg13g2_inv_4 U3201 (.A(n3061), .Y(n3055));
sg13g2_o21ai_1 U3202 (.A1(n4327), .A2(n3059), .B1(n3063), .Y(n3061));
sg13g2_a21oi_2 U3203 (.A1(data_i_26_), .A2(n4307), .B1(n3064), .Y(n3063));
sg13g2_nor2_2 U3204 (.A(n555), .B(n721), .Y(n3064));
sg13g2_inv_4 U3205 (.A(mixcol_data_o_26), .Y(n721));
sg13g2_inv_4 U3206 (.A(subbytes_data_o_26), .Y(n3059));
sg13g2_a21oi_2 U3208 (.A1(n2244), .A2(n3067), .B1(n3068), .Y(n3066));
sg13g2_nor2_2 U3209 (.A(n3069), .B(n2248), .Y(n3068));
sg13g2_o21ai_1 U3210 (.A1(n4167), .A2(n3069), .B1(n3070), .Y(n3067));
sg13g2_a21oi_2 U3211 (.A1(n4315), .A2(n3071), .B1(n3072), .Y(n3070));
sg13g2_nor2_2 U3212 (.A(n4164), .B(n723), .Y(n3072));
sg13g2_inv_4 U3213 (.A(n3071), .Y(n3065));
sg13g2_o21ai_1 U3214 (.A1(n4325), .A2(n3069), .B1(n3073), .Y(n3071));
sg13g2_a21oi_2 U3215 (.A1(data_i_25_), .A2(n4307), .B1(n3074), .Y(n3073));
sg13g2_nor2_2 U3216 (.A(n555), .B(n723), .Y(n3074));
sg13g2_inv_4 U3217 (.A(mixcol_data_o_25), .Y(n723));
sg13g2_inv_4 U3218 (.A(subbytes_data_o_25), .Y(n3069));
sg13g2_a21oi_2 U3220 (.A1(n4313), .A2(n3077), .B1(n3078), .Y(n3076));
sg13g2_nor2_2 U3221 (.A(n3079), .B(n2248), .Y(n3078));
sg13g2_o21ai_1 U3222 (.A1(n4167), .A2(n3079), .B1(n3080), .Y(n3077));
sg13g2_a21oi_2 U3223 (.A1(n4315), .A2(n3081), .B1(n3082), .Y(n3080));
sg13g2_nor2_2 U3224 (.A(n4165), .B(n725), .Y(n3082));
sg13g2_inv_4 U3225 (.A(n3081), .Y(n3075));
sg13g2_o21ai_1 U3226 (.A1(n4329), .A2(n3079), .B1(n3083), .Y(n3081));
sg13g2_a21oi_2 U3227 (.A1(data_i_24_), .A2(n4307), .B1(n3084), .Y(n3083));
sg13g2_nor2_2 U3228 (.A(n555), .B(n725), .Y(n3084));
sg13g2_inv_4 U3229 (.A(mixcol_data_o_24), .Y(n725));
sg13g2_inv_4 U3230 (.A(subbytes_data_o_24), .Y(n3079));
sg13g2_a21oi_2 U3232 (.A1(n4313), .A2(n3087), .B1(n3088), .Y(n3086));
sg13g2_nor2_2 U3233 (.A(n3089), .B(n2248), .Y(n3088));
sg13g2_o21ai_1 U3234 (.A1(n553), .A2(n3089), .B1(n3090), .Y(n3087));
sg13g2_a21oi_2 U3235 (.A1(n4315), .A2(n3091), .B1(n3092), .Y(n3090));
sg13g2_nor2_2 U3236 (.A(n4165), .B(n727), .Y(n3092));
sg13g2_inv_4 U3237 (.A(n3091), .Y(n3085));
sg13g2_o21ai_1 U3238 (.A1(n4325), .A2(n3089), .B1(n3093), .Y(n3091));
sg13g2_a21oi_2 U3239 (.A1(data_i_23_), .A2(n4307), .B1(n3094), .Y(n3093));
sg13g2_nor2_2 U3240 (.A(n555), .B(n727), .Y(n3094));
sg13g2_inv_4 U3241 (.A(mixcol_data_o_23), .Y(n727));
sg13g2_inv_4 U3242 (.A(subbytes_data_o_23), .Y(n3089));
sg13g2_a21oi_2 U3244 (.A1(n4313), .A2(n3097), .B1(n3098), .Y(n3096));
sg13g2_nor2_2 U3245 (.A(n3099), .B(n2248), .Y(n3098));
sg13g2_o21ai_1 U3246 (.A1(n553), .A2(n3099), .B1(n3100), .Y(n3097));
sg13g2_a21oi_2 U3247 (.A1(n4315), .A2(n3101), .B1(n3102), .Y(n3100));
sg13g2_nor2_2 U3248 (.A(n4164), .B(n729), .Y(n3102));
sg13g2_inv_4 U3249 (.A(n3101), .Y(n3095));
sg13g2_o21ai_1 U3250 (.A1(n4330), .A2(n3099), .B1(n3103), .Y(n3101));
sg13g2_a21oi_2 U3251 (.A1(data_i_22_), .A2(n4307), .B1(n3104), .Y(n3103));
sg13g2_nor2_2 U3252 (.A(n555), .B(n729), .Y(n3104));
sg13g2_inv_4 U3253 (.A(mixcol_data_o_22), .Y(n729));
sg13g2_inv_4 U3254 (.A(subbytes_data_o_22), .Y(n3099));
sg13g2_a21oi_2 U3256 (.A1(n2244), .A2(n3107), .B1(n3108), .Y(n3106));
sg13g2_nor2_2 U3257 (.A(n3109), .B(n2248), .Y(n3108));
sg13g2_o21ai_1 U3258 (.A1(n553), .A2(n3109), .B1(n3110), .Y(n3107));
sg13g2_a21oi_2 U3259 (.A1(n4315), .A2(n3111), .B1(n3112), .Y(n3110));
sg13g2_nor2_2 U3260 (.A(n4165), .B(n731), .Y(n3112));
sg13g2_inv_4 U3261 (.A(n3111), .Y(n3105));
sg13g2_o21ai_1 U3262 (.A1(n4326), .A2(n3109), .B1(n3113), .Y(n3111));
sg13g2_a21oi_2 U3263 (.A1(data_i_21_), .A2(n4307), .B1(n3114), .Y(n3113));
sg13g2_nor2_2 U3264 (.A(n555), .B(n731), .Y(n3114));
sg13g2_inv_4 U3265 (.A(mixcol_data_o_21), .Y(n731));
sg13g2_inv_4 U3266 (.A(subbytes_data_o_21), .Y(n3109));
sg13g2_a21oi_2 U3268 (.A1(n4312), .A2(n3117), .B1(n3118), .Y(n3116));
sg13g2_nor2_2 U3269 (.A(n3119), .B(n2248), .Y(n3118));
sg13g2_o21ai_1 U3270 (.A1(n553), .A2(n3119), .B1(n3120), .Y(n3117));
sg13g2_a21oi_2 U3271 (.A1(n4315), .A2(n3121), .B1(n3122), .Y(n3120));
sg13g2_nor2_2 U3272 (.A(n4165), .B(n733), .Y(n3122));
sg13g2_inv_4 U3273 (.A(n3121), .Y(n3115));
sg13g2_o21ai_1 U3274 (.A1(n4330), .A2(n3119), .B1(n3123), .Y(n3121));
sg13g2_a21oi_2 U3275 (.A1(data_i_20_), .A2(n4307), .B1(n3124), .Y(n3123));
sg13g2_nor2_2 U3276 (.A(n555), .B(n733), .Y(n3124));
sg13g2_inv_4 U3277 (.A(mixcol_data_o_20), .Y(n733));
sg13g2_inv_4 U3278 (.A(subbytes_data_o_20), .Y(n3119));
sg13g2_a21oi_2 U3280 (.A1(n2244), .A2(n3127), .B1(n3128), .Y(n3126));
sg13g2_nor2_2 U3281 (.A(n3129), .B(n2248), .Y(n3128));
sg13g2_o21ai_1 U3282 (.A1(n4167), .A2(n3129), .B1(n3130), .Y(n3127));
sg13g2_a21oi_2 U3283 (.A1(n4315), .A2(n3131), .B1(n3132), .Y(n3130));
sg13g2_nor2_2 U3284 (.A(n4165), .B(n735), .Y(n3132));
sg13g2_inv_4 U3285 (.A(n3131), .Y(n3125));
sg13g2_o21ai_1 U3286 (.A1(n4330), .A2(n3129), .B1(n3133), .Y(n3131));
sg13g2_a21oi_2 U3287 (.A1(data_i_1_), .A2(n4307), .B1(n3134), .Y(n3133));
sg13g2_nor2_2 U3288 (.A(n555), .B(n735), .Y(n3134));
sg13g2_inv_4 U3289 (.A(mixcol_data_o_1), .Y(n735));
sg13g2_inv_4 U3290 (.A(subbytes_data_o_1), .Y(n3129));
sg13g2_a21oi_2 U3292 (.A1(n2244), .A2(n3137), .B1(n3138), .Y(n3136));
sg13g2_nor2_2 U3293 (.A(n3139), .B(n2248), .Y(n3138));
sg13g2_o21ai_1 U3294 (.A1(n553), .A2(n3139), .B1(n3140), .Y(n3137));
sg13g2_a21oi_2 U3295 (.A1(n4315), .A2(n3141), .B1(n3142), .Y(n3140));
sg13g2_nor2_2 U3296 (.A(n4165), .B(n737), .Y(n3142));
sg13g2_inv_4 U3297 (.A(n3141), .Y(n3135));
sg13g2_o21ai_1 U3298 (.A1(n4325), .A2(n3139), .B1(n3143), .Y(n3141));
sg13g2_a21oi_2 U3299 (.A1(data_i_19_), .A2(n4308), .B1(n3144), .Y(n3143));
sg13g2_nor2_2 U3300 (.A(n555), .B(n737), .Y(n3144));
sg13g2_inv_4 U3301 (.A(mixcol_data_o_19), .Y(n737));
sg13g2_inv_4 U3302 (.A(subbytes_data_o_19), .Y(n3139));
sg13g2_o21ai_1 U3303 (.A1(n4332), .A2(n3145), .B1(n3146), .Y(addroundkey_data_i_18));
sg13g2_a21oi_2 U3304 (.A1(n4313), .A2(n3147), .B1(n3148), .Y(n3146));
sg13g2_nor2_2 U3305 (.A(n3149), .B(n4310), .Y(n3148));
sg13g2_o21ai_1 U3306 (.A1(n4167), .A2(n3149), .B1(n3150), .Y(n3147));
sg13g2_a21oi_2 U3307 (.A1(n4315), .A2(n3151), .B1(n3152), .Y(n3150));
sg13g2_nor2_2 U3308 (.A(n4165), .B(n739), .Y(n3152));
sg13g2_inv_4 U3309 (.A(n3151), .Y(n3145));
sg13g2_o21ai_1 U3310 (.A1(n4326), .A2(n3149), .B1(n3153), .Y(n3151));
sg13g2_a21oi_2 U3311 (.A1(data_i_18_), .A2(n4308), .B1(n3154), .Y(n3153));
sg13g2_nor2_2 U3312 (.A(n555), .B(n739), .Y(n3154));
sg13g2_inv_4 U3313 (.A(mixcol_data_o_18), .Y(n739));
sg13g2_inv_4 U3314 (.A(subbytes_data_o_18), .Y(n3149));
sg13g2_a21oi_2 U3316 (.A1(n4313), .A2(n3157), .B1(n3158), .Y(n3156));
sg13g2_nor2_2 U3317 (.A(n3159), .B(n2248), .Y(n3158));
sg13g2_o21ai_1 U3318 (.A1(n553), .A2(n3159), .B1(n3160), .Y(n3157));
sg13g2_a21oi_2 U3319 (.A1(n4315), .A2(n3161), .B1(n3162), .Y(n3160));
sg13g2_nor2_2 U3320 (.A(n4164), .B(n741), .Y(n3162));
sg13g2_inv_4 U3321 (.A(n3161), .Y(n3155));
sg13g2_o21ai_1 U3322 (.A1(n4328), .A2(n3159), .B1(n3163), .Y(n3161));
sg13g2_a21oi_2 U3323 (.A1(data_i_17_), .A2(n4307), .B1(n3164), .Y(n3163));
sg13g2_nor2_2 U3324 (.A(n555), .B(n741), .Y(n3164));
sg13g2_inv_4 U3325 (.A(mixcol_data_o_17), .Y(n741));
sg13g2_inv_4 U3326 (.A(subbytes_data_o_17), .Y(n3159));
sg13g2_a21oi_2 U3328 (.A1(n4313), .A2(n3167), .B1(n3168), .Y(n3166));
sg13g2_nor2_2 U3329 (.A(n3169), .B(n2248), .Y(n3168));
sg13g2_o21ai_1 U3330 (.A1(n4167), .A2(n3169), .B1(n3170), .Y(n3167));
sg13g2_a21oi_2 U3331 (.A1(n4315), .A2(n3171), .B1(n3172), .Y(n3170));
sg13g2_nor2_2 U3332 (.A(n4165), .B(n743), .Y(n3172));
sg13g2_inv_4 U3333 (.A(n3171), .Y(n3165));
sg13g2_o21ai_1 U3334 (.A1(n4326), .A2(n3169), .B1(n3173), .Y(n3171));
sg13g2_a21oi_2 U3335 (.A1(data_i_16_), .A2(n4308), .B1(n3174), .Y(n3173));
sg13g2_nor2_2 U3336 (.A(n555), .B(n743), .Y(n3174));
sg13g2_inv_4 U3337 (.A(mixcol_data_o_16), .Y(n743));
sg13g2_inv_4 U3338 (.A(subbytes_data_o_16), .Y(n3169));
sg13g2_a21oi_2 U3340 (.A1(n2244), .A2(n3177), .B1(n3178), .Y(n3176));
sg13g2_nor2_2 U3341 (.A(n3179), .B(n2248), .Y(n3178));
sg13g2_o21ai_1 U3342 (.A1(n4167), .A2(n3179), .B1(n3180), .Y(n3177));
sg13g2_a21oi_2 U3343 (.A1(n4315), .A2(n3181), .B1(n3182), .Y(n3180));
sg13g2_nor2_2 U3344 (.A(n4165), .B(n745), .Y(n3182));
sg13g2_inv_4 U3345 (.A(n3181), .Y(n3175));
sg13g2_o21ai_1 U3346 (.A1(n4325), .A2(n3179), .B1(n3183), .Y(n3181));
sg13g2_a21oi_2 U3347 (.A1(data_i_15_), .A2(n4307), .B1(n3184), .Y(n3183));
sg13g2_nor2_2 U3348 (.A(n555), .B(n745), .Y(n3184));
sg13g2_inv_4 U3349 (.A(mixcol_data_o_15), .Y(n745));
sg13g2_inv_4 U3350 (.A(subbytes_data_o_15), .Y(n3179));
sg13g2_a21oi_2 U3352 (.A1(n2244), .A2(n3187), .B1(n3188), .Y(n3186));
sg13g2_nor2_2 U3353 (.A(n3189), .B(n2248), .Y(n3188));
sg13g2_o21ai_1 U3354 (.A1(n553), .A2(n3189), .B1(n3190), .Y(n3187));
sg13g2_a21oi_2 U3355 (.A1(n4315), .A2(n3191), .B1(n3192), .Y(n3190));
sg13g2_nor2_2 U3356 (.A(n4165), .B(n747), .Y(n3192));
sg13g2_inv_4 U3357 (.A(n3191), .Y(n3185));
sg13g2_o21ai_1 U3358 (.A1(n4329), .A2(n3189), .B1(n3193), .Y(n3191));
sg13g2_a21oi_2 U3359 (.A1(data_i_14_), .A2(n4307), .B1(n3194), .Y(n3193));
sg13g2_nor2_2 U3360 (.A(n555), .B(n747), .Y(n3194));
sg13g2_inv_4 U3361 (.A(mixcol_data_o_14), .Y(n747));
sg13g2_inv_4 U3362 (.A(subbytes_data_o_14), .Y(n3189));
sg13g2_a21oi_2 U3364 (.A1(n2244), .A2(n3197), .B1(n3198), .Y(n3196));
sg13g2_nor2_2 U3365 (.A(n3199), .B(n2248), .Y(n3198));
sg13g2_o21ai_1 U3366 (.A1(n553), .A2(n3199), .B1(n3200), .Y(n3197));
sg13g2_a21oi_2 U3367 (.A1(n4315), .A2(n3201), .B1(n3202), .Y(n3200));
sg13g2_nor2_2 U3368 (.A(n4164), .B(n749), .Y(n3202));
sg13g2_inv_4 U3369 (.A(n3201), .Y(n3195));
sg13g2_o21ai_1 U3370 (.A1(n4326), .A2(n3199), .B1(n3203), .Y(n3201));
sg13g2_a21oi_2 U3371 (.A1(data_i_13_), .A2(n4308), .B1(n3204), .Y(n3203));
sg13g2_nor2_2 U3372 (.A(n555), .B(n749), .Y(n3204));
sg13g2_inv_4 U3373 (.A(mixcol_data_o_13), .Y(n749));
sg13g2_inv_4 U3374 (.A(subbytes_data_o_13), .Y(n3199));
sg13g2_nor2_2 U3377 (.A(n3209), .B(n2248), .Y(n3208));
sg13g2_o21ai_1 U3378 (.A1(n553), .A2(n3209), .B1(n3210), .Y(n3207));
sg13g2_a21oi_2 U3379 (.A1(n4315), .A2(n3211), .B1(n3212), .Y(n3210));
sg13g2_nor2_2 U3380 (.A(n4164), .B(n751), .Y(n3212));
sg13g2_inv_4 U3381 (.A(n3211), .Y(n3205));
sg13g2_o21ai_1 U3382 (.A1(n4330), .A2(n3209), .B1(n3213), .Y(n3211));
sg13g2_a21oi_2 U3383 (.A1(data_i_12_), .A2(n2253), .B1(n3214), .Y(n3213));
sg13g2_nor2_2 U3384 (.A(n555), .B(n751), .Y(n3214));
sg13g2_inv_4 U3385 (.A(mixcol_data_o_12), .Y(n751));
sg13g2_inv_4 U3386 (.A(subbytes_data_o_12), .Y(n3209));
sg13g2_a21oi_2 U3388 (.A1(n4313), .A2(n3217), .B1(n3218), .Y(n3216));
sg13g2_nor2_2 U3389 (.A(n3219), .B(n2248), .Y(n3218));
sg13g2_o21ai_1 U3390 (.A1(n4167), .A2(n3219), .B1(n3220), .Y(n3217));
sg13g2_a21oi_2 U3391 (.A1(n4315), .A2(n3221), .B1(n3222), .Y(n3220));
sg13g2_nor2_2 U3392 (.A(n4165), .B(n753), .Y(n3222));
sg13g2_inv_4 U3393 (.A(n3221), .Y(n3215));
sg13g2_o21ai_1 U3394 (.A1(n4325), .A2(n3219), .B1(n3223), .Y(n3221));
sg13g2_a21oi_2 U3395 (.A1(data_i_127_), .A2(n4308), .B1(n3224), .Y(n3223));
sg13g2_nor2_2 U3396 (.A(n555), .B(n753), .Y(n3224));
sg13g2_inv_4 U3397 (.A(mixcol_data_o_127), .Y(n753));
sg13g2_inv_4 U3398 (.A(subbytes_data_o_127), .Y(n3219));
sg13g2_a21oi_2 U3400 (.A1(n2244), .A2(n3227), .B1(n3228), .Y(n3226));
sg13g2_nor2_2 U3401 (.A(n3229), .B(n2248), .Y(n3228));
sg13g2_o21ai_1 U3402 (.A1(n4167), .A2(n3229), .B1(n3230), .Y(n3227));
sg13g2_a21oi_2 U3403 (.A1(n4315), .A2(n3231), .B1(n3232), .Y(n3230));
sg13g2_nor2_2 U3404 (.A(n4164), .B(n755), .Y(n3232));
sg13g2_inv_4 U3405 (.A(n3231), .Y(n3225));
sg13g2_o21ai_1 U3406 (.A1(n4327), .A2(n3229), .B1(n3233), .Y(n3231));
sg13g2_a21oi_2 U3407 (.A1(data_i_126_), .A2(n4307), .B1(n3234), .Y(n3233));
sg13g2_nor2_2 U3408 (.A(n555), .B(n755), .Y(n3234));
sg13g2_inv_4 U3409 (.A(mixcol_data_o_126), .Y(n755));
sg13g2_inv_4 U3410 (.A(subbytes_data_o_126), .Y(n3229));
sg13g2_a21oi_2 U3412 (.A1(n4313), .A2(n3237), .B1(n3238), .Y(n3236));
sg13g2_nor2_2 U3413 (.A(n3239), .B(n2248), .Y(n3238));
sg13g2_o21ai_1 U3414 (.A1(n553), .A2(n3239), .B1(n3240), .Y(n3237));
sg13g2_a21oi_2 U3415 (.A1(n4315), .A2(n3241), .B1(n3242), .Y(n3240));
sg13g2_nor2_2 U3416 (.A(n4165), .B(n757), .Y(n3242));
sg13g2_inv_4 U3417 (.A(n3241), .Y(n3235));
sg13g2_o21ai_1 U3418 (.A1(n4327), .A2(n3239), .B1(n3243), .Y(n3241));
sg13g2_a21oi_2 U3419 (.A1(data_i_125_), .A2(n4308), .B1(n3244), .Y(n3243));
sg13g2_nor2_2 U3420 (.A(n555), .B(n757), .Y(n3244));
sg13g2_inv_4 U3421 (.A(mixcol_data_o_125), .Y(n757));
sg13g2_inv_4 U3422 (.A(subbytes_data_o_125), .Y(n3239));
sg13g2_a21oi_2 U3424 (.A1(n4313), .A2(n3247), .B1(n3248), .Y(n3246));
sg13g2_nor2_2 U3425 (.A(n3249), .B(n2248), .Y(n3248));
sg13g2_o21ai_1 U3426 (.A1(n4167), .A2(n3249), .B1(n3250), .Y(n3247));
sg13g2_a21oi_2 U3427 (.A1(n4315), .A2(n3251), .B1(n3252), .Y(n3250));
sg13g2_nor2_2 U3428 (.A(n4164), .B(n759), .Y(n3252));
sg13g2_inv_4 U3429 (.A(n3251), .Y(n3245));
sg13g2_o21ai_1 U3430 (.A1(n4327), .A2(n3249), .B1(n3253), .Y(n3251));
sg13g2_a21oi_2 U3431 (.A1(data_i_124_), .A2(n4308), .B1(n3254), .Y(n3253));
sg13g2_nor2_2 U3432 (.A(n555), .B(n759), .Y(n3254));
sg13g2_inv_4 U3433 (.A(mixcol_data_o_124), .Y(n759));
sg13g2_inv_4 U3434 (.A(subbytes_data_o_124), .Y(n3249));
sg13g2_nor2_2 U3437 (.A(n3259), .B(n2248), .Y(n3258));
sg13g2_o21ai_1 U3438 (.A1(n4167), .A2(n3259), .B1(n3260), .Y(n3257));
sg13g2_a21oi_2 U3439 (.A1(n4315), .A2(n3261), .B1(n3262), .Y(n3260));
sg13g2_nor2_2 U3440 (.A(n4165), .B(n761), .Y(n3262));
sg13g2_inv_4 U3441 (.A(n3261), .Y(n3255));
sg13g2_o21ai_1 U3442 (.A1(n4326), .A2(n3259), .B1(n3263), .Y(n3261));
sg13g2_a21oi_2 U3443 (.A1(data_i_123_), .A2(n4308), .B1(n3264), .Y(n3263));
sg13g2_nor2_2 U3444 (.A(n555), .B(n761), .Y(n3264));
sg13g2_inv_4 U3445 (.A(mixcol_data_o_123), .Y(n761));
sg13g2_inv_4 U3446 (.A(subbytes_data_o_123), .Y(n3259));
sg13g2_nor2_2 U3449 (.A(n3269), .B(n2248), .Y(n3268));
sg13g2_o21ai_1 U3450 (.A1(n553), .A2(n3269), .B1(n3270), .Y(n3267));
sg13g2_a21oi_2 U3451 (.A1(n4315), .A2(n3271), .B1(n3272), .Y(n3270));
sg13g2_nor2_2 U3452 (.A(n4165), .B(n763), .Y(n3272));
sg13g2_inv_4 U3453 (.A(n3271), .Y(n3265));
sg13g2_o21ai_1 U3454 (.A1(n4328), .A2(n3269), .B1(n3273), .Y(n3271));
sg13g2_a21oi_2 U3455 (.A1(data_i_122_), .A2(n4308), .B1(n3274), .Y(n3273));
sg13g2_nor2_2 U3456 (.A(n555), .B(n763), .Y(n3274));
sg13g2_inv_4 U3457 (.A(mixcol_data_o_122), .Y(n763));
sg13g2_inv_4 U3458 (.A(subbytes_data_o_122), .Y(n3269));
sg13g2_nor2_2 U3461 (.A(n3279), .B(n2248), .Y(n3278));
sg13g2_o21ai_1 U3462 (.A1(n4167), .A2(n3279), .B1(n3280), .Y(n3277));
sg13g2_a21oi_2 U3463 (.A1(n4315), .A2(n3281), .B1(n3282), .Y(n3280));
sg13g2_nor2_2 U3464 (.A(n4165), .B(n765), .Y(n3282));
sg13g2_inv_4 U3465 (.A(n3281), .Y(n3275));
sg13g2_o21ai_1 U3466 (.A1(n4327), .A2(n3279), .B1(n3283), .Y(n3281));
sg13g2_a21oi_2 U3467 (.A1(data_i_121_), .A2(n2253), .B1(n3284), .Y(n3283));
sg13g2_nor2_2 U3468 (.A(n555), .B(n765), .Y(n3284));
sg13g2_inv_4 U3469 (.A(mixcol_data_o_121), .Y(n765));
sg13g2_inv_4 U3470 (.A(subbytes_data_o_121), .Y(n3279));
sg13g2_nor2_2 U3473 (.A(n3289), .B(n2248), .Y(n3288));
sg13g2_o21ai_1 U3474 (.A1(n553), .A2(n3289), .B1(n3290), .Y(n3287));
sg13g2_a21oi_2 U3475 (.A1(n4315), .A2(n3291), .B1(n3292), .Y(n3290));
sg13g2_nor2_2 U3476 (.A(n4164), .B(n767), .Y(n3292));
sg13g2_inv_4 U3477 (.A(n3291), .Y(n3285));
sg13g2_o21ai_1 U3478 (.A1(n4330), .A2(n3289), .B1(n3293), .Y(n3291));
sg13g2_a21oi_2 U3479 (.A1(data_i_120_), .A2(n2253), .B1(n3294), .Y(n3293));
sg13g2_nor2_2 U3480 (.A(n555), .B(n767), .Y(n3294));
sg13g2_inv_4 U3481 (.A(mixcol_data_o_120), .Y(n767));
sg13g2_inv_4 U3482 (.A(subbytes_data_o_120), .Y(n3289));
sg13g2_nor2_2 U3485 (.A(n3299), .B(n2248), .Y(n3298));
sg13g2_o21ai_1 U3486 (.A1(n4167), .A2(n3299), .B1(n3300), .Y(n3297));
sg13g2_a21oi_2 U3487 (.A1(n4315), .A2(n3301), .B1(n3302), .Y(n3300));
sg13g2_nor2_2 U3488 (.A(n4164), .B(n769), .Y(n3302));
sg13g2_inv_4 U3489 (.A(n3301), .Y(n3295));
sg13g2_o21ai_1 U3490 (.A1(n4328), .A2(n3299), .B1(n3303), .Y(n3301));
sg13g2_a21oi_2 U3491 (.A1(data_i_11_), .A2(n4308), .B1(n3304), .Y(n3303));
sg13g2_nor2_2 U3492 (.A(n555), .B(n769), .Y(n3304));
sg13g2_inv_4 U3493 (.A(mixcol_data_o_11), .Y(n769));
sg13g2_inv_4 U3494 (.A(subbytes_data_o_11), .Y(n3299));
sg13g2_nor2_2 U3497 (.A(n3309), .B(n2248), .Y(n3308));
sg13g2_o21ai_1 U3498 (.A1(n553), .A2(n3309), .B1(n3310), .Y(n3307));
sg13g2_a21oi_2 U3499 (.A1(n4315), .A2(n3311), .B1(n3312), .Y(n3310));
sg13g2_nor2_2 U3500 (.A(n4164), .B(n771), .Y(n3312));
sg13g2_inv_4 U3501 (.A(n3311), .Y(n3305));
sg13g2_o21ai_1 U3502 (.A1(n4328), .A2(n3309), .B1(n3313), .Y(n3311));
sg13g2_a21oi_2 U3503 (.A1(data_i_119_), .A2(n2253), .B1(n3314), .Y(n3313));
sg13g2_nor2_2 U3504 (.A(n555), .B(n771), .Y(n3314));
sg13g2_inv_4 U3505 (.A(mixcol_data_o_119), .Y(n771));
sg13g2_inv_4 U3506 (.A(subbytes_data_o_119), .Y(n3309));
sg13g2_nor2_2 U3509 (.A(n3319), .B(n2248), .Y(n3318));
sg13g2_o21ai_1 U3510 (.A1(n4167), .A2(n3319), .B1(n3320), .Y(n3317));
sg13g2_a21oi_2 U3511 (.A1(n4315), .A2(n3321), .B1(n3322), .Y(n3320));
sg13g2_nor2_2 U3512 (.A(n4164), .B(n773), .Y(n3322));
sg13g2_inv_4 U3513 (.A(n3321), .Y(n3315));
sg13g2_o21ai_1 U3514 (.A1(n4329), .A2(n3319), .B1(n3323), .Y(n3321));
sg13g2_a21oi_2 U3515 (.A1(data_i_118_), .A2(n4308), .B1(n3324), .Y(n3323));
sg13g2_nor2_2 U3516 (.A(n555), .B(n773), .Y(n3324));
sg13g2_inv_4 U3517 (.A(mixcol_data_o_118), .Y(n773));
sg13g2_inv_4 U3518 (.A(subbytes_data_o_118), .Y(n3319));
sg13g2_nor2_2 U3521 (.A(n3329), .B(n2248), .Y(n3328));
sg13g2_o21ai_1 U3522 (.A1(n553), .A2(n3329), .B1(n3330), .Y(n3327));
sg13g2_a21oi_2 U3523 (.A1(n4315), .A2(n3331), .B1(n3332), .Y(n3330));
sg13g2_nor2_2 U3524 (.A(n4164), .B(n775), .Y(n3332));
sg13g2_inv_4 U3525 (.A(n3331), .Y(n3325));
sg13g2_o21ai_1 U3526 (.A1(n4329), .A2(n3329), .B1(n3333), .Y(n3331));
sg13g2_a21oi_2 U3527 (.A1(data_i_117_), .A2(n4307), .B1(n3334), .Y(n3333));
sg13g2_nor2_2 U3528 (.A(n555), .B(n775), .Y(n3334));
sg13g2_inv_4 U3529 (.A(mixcol_data_o_117), .Y(n775));
sg13g2_inv_4 U3530 (.A(subbytes_data_o_117), .Y(n3329));
sg13g2_nor2_2 U3533 (.A(n3339), .B(n2248), .Y(n3338));
sg13g2_o21ai_1 U3534 (.A1(n4167), .A2(n3339), .B1(n3340), .Y(n3337));
sg13g2_a21oi_2 U3535 (.A1(n4315), .A2(n3341), .B1(n3342), .Y(n3340));
sg13g2_nor2_2 U3536 (.A(n4164), .B(n777), .Y(n3342));
sg13g2_inv_4 U3537 (.A(n3341), .Y(n3335));
sg13g2_o21ai_1 U3538 (.A1(n4329), .A2(n3339), .B1(n3343), .Y(n3341));
sg13g2_a21oi_2 U3539 (.A1(data_i_116_), .A2(n4307), .B1(n3344), .Y(n3343));
sg13g2_nor2_2 U3540 (.A(n555), .B(n777), .Y(n3344));
sg13g2_inv_4 U3541 (.A(mixcol_data_o_116), .Y(n777));
sg13g2_inv_4 U3542 (.A(subbytes_data_o_116), .Y(n3339));
sg13g2_o21ai_1 U3543 (.A1(n4332), .A2(n3345), .B1(n3346), .Y(addroundkey_data_i_115));
sg13g2_nor2_2 U3545 (.A(n3349), .B(n2248), .Y(n3348));
sg13g2_o21ai_1 U3546 (.A1(n4167), .A2(n3349), .B1(n3350), .Y(n3347));
sg13g2_a21oi_2 U3547 (.A1(n4315), .A2(n3351), .B1(n3352), .Y(n3350));
sg13g2_nor2_2 U3548 (.A(n4165), .B(n779), .Y(n3352));
sg13g2_inv_4 U3549 (.A(n3351), .Y(n3345));
sg13g2_o21ai_1 U3550 (.A1(n4326), .A2(n3349), .B1(n3353), .Y(n3351));
sg13g2_a21oi_2 U3551 (.A1(data_i_115_), .A2(n4307), .B1(n3354), .Y(n3353));
sg13g2_nor2_2 U3552 (.A(n555), .B(n779), .Y(n3354));
sg13g2_inv_4 U3553 (.A(mixcol_data_o_115), .Y(n779));
sg13g2_inv_4 U3554 (.A(subbytes_data_o_115), .Y(n3349));
sg13g2_nor2_2 U3557 (.A(n3359), .B(n2248), .Y(n3358));
sg13g2_o21ai_1 U3558 (.A1(n553), .A2(n3359), .B1(n3360), .Y(n3357));
sg13g2_a21oi_2 U3559 (.A1(n4315), .A2(n3361), .B1(n3362), .Y(n3360));
sg13g2_nor2_2 U3560 (.A(n4164), .B(n781), .Y(n3362));
sg13g2_inv_4 U3561 (.A(n3361), .Y(n3355));
sg13g2_o21ai_1 U3562 (.A1(n4328), .A2(n3359), .B1(n3363), .Y(n3361));
sg13g2_a21oi_2 U3563 (.A1(data_i_114_), .A2(n4307), .B1(n3364), .Y(n3363));
sg13g2_nor2_2 U3564 (.A(n555), .B(n781), .Y(n3364));
sg13g2_inv_4 U3565 (.A(mixcol_data_o_114), .Y(n781));
sg13g2_inv_4 U3566 (.A(subbytes_data_o_114), .Y(n3359));
sg13g2_o21ai_1 U3567 (.A1(n4332), .A2(n3365), .B1(n3366), .Y(addroundkey_data_i_113));
sg13g2_nor2_2 U3569 (.A(n3369), .B(n2248), .Y(n3368));
sg13g2_o21ai_1 U3570 (.A1(n4167), .A2(n3369), .B1(n3370), .Y(n3367));
sg13g2_a21oi_2 U3571 (.A1(n4315), .A2(n3371), .B1(n3372), .Y(n3370));
sg13g2_nor2_2 U3572 (.A(n4165), .B(n783), .Y(n3372));
sg13g2_inv_4 U3573 (.A(n3371), .Y(n3365));
sg13g2_o21ai_1 U3574 (.A1(n4325), .A2(n3369), .B1(n3373), .Y(n3371));
sg13g2_a21oi_2 U3575 (.A1(data_i_113_), .A2(n4307), .B1(n3374), .Y(n3373));
sg13g2_nor2_2 U3576 (.A(n555), .B(n783), .Y(n3374));
sg13g2_inv_4 U3577 (.A(mixcol_data_o_113), .Y(n783));
sg13g2_inv_4 U3578 (.A(subbytes_data_o_113), .Y(n3369));
sg13g2_nor2_2 U3581 (.A(n3379), .B(n2248), .Y(n3378));
sg13g2_o21ai_1 U3582 (.A1(n553), .A2(n3379), .B1(n3380), .Y(n3377));
sg13g2_a21oi_2 U3583 (.A1(n4315), .A2(n3381), .B1(n3382), .Y(n3380));
sg13g2_nor2_2 U3584 (.A(n4165), .B(n785), .Y(n3382));
sg13g2_inv_4 U3585 (.A(n3381), .Y(n3375));
sg13g2_o21ai_1 U3586 (.A1(n4328), .A2(n3379), .B1(n3383), .Y(n3381));
sg13g2_a21oi_2 U3587 (.A1(data_i_112_), .A2(n4307), .B1(n3384), .Y(n3383));
sg13g2_nor2_2 U3588 (.A(n555), .B(n785), .Y(n3384));
sg13g2_inv_4 U3589 (.A(mixcol_data_o_112), .Y(n785));
sg13g2_inv_4 U3590 (.A(subbytes_data_o_112), .Y(n3379));
sg13g2_o21ai_1 U3591 (.A1(n4332), .A2(n3385), .B1(n3386), .Y(addroundkey_data_i_111));
sg13g2_nor2_2 U3593 (.A(n3389), .B(n2248), .Y(n3388));
sg13g2_o21ai_1 U3594 (.A1(n4167), .A2(n3389), .B1(n3390), .Y(n3387));
sg13g2_a21oi_2 U3595 (.A1(n4315), .A2(n3391), .B1(n3392), .Y(n3390));
sg13g2_nor2_2 U3596 (.A(n4165), .B(n787), .Y(n3392));
sg13g2_inv_4 U3597 (.A(n3391), .Y(n3385));
sg13g2_o21ai_1 U3598 (.A1(n4326), .A2(n3389), .B1(n3393), .Y(n3391));
sg13g2_a21oi_2 U3599 (.A1(data_i_111_), .A2(n4307), .B1(n3394), .Y(n3393));
sg13g2_nor2_2 U3600 (.A(n555), .B(n787), .Y(n3394));
sg13g2_inv_4 U3601 (.A(mixcol_data_o_111), .Y(n787));
sg13g2_inv_4 U3602 (.A(subbytes_data_o_111), .Y(n3389));
sg13g2_nor2_2 U3605 (.A(n3399), .B(n2248), .Y(n3398));
sg13g2_o21ai_1 U3606 (.A1(n4167), .A2(n3399), .B1(n3400), .Y(n3397));
sg13g2_a21oi_2 U3607 (.A1(n4315), .A2(n3401), .B1(n3402), .Y(n3400));
sg13g2_nor2_2 U3608 (.A(n4165), .B(n789), .Y(n3402));
sg13g2_inv_4 U3609 (.A(n3401), .Y(n3395));
sg13g2_o21ai_1 U3610 (.A1(n4328), .A2(n3399), .B1(n3403), .Y(n3401));
sg13g2_a21oi_2 U3611 (.A1(data_i_110_), .A2(n4307), .B1(n3404), .Y(n3403));
sg13g2_nor2_2 U3612 (.A(n555), .B(n789), .Y(n3404));
sg13g2_inv_4 U3613 (.A(mixcol_data_o_110), .Y(n789));
sg13g2_inv_4 U3614 (.A(subbytes_data_o_110), .Y(n3399));
sg13g2_nor2_2 U3617 (.A(n3409), .B(n2248), .Y(n3408));
sg13g2_o21ai_1 U3618 (.A1(n553), .A2(n3409), .B1(n3410), .Y(n3407));
sg13g2_a21oi_2 U3619 (.A1(n4315), .A2(n3411), .B1(n3412), .Y(n3410));
sg13g2_nor2_2 U3620 (.A(n4165), .B(n791), .Y(n3412));
sg13g2_inv_4 U3621 (.A(n3411), .Y(n3405));
sg13g2_o21ai_1 U3622 (.A1(n4326), .A2(n3409), .B1(n3413), .Y(n3411));
sg13g2_a21oi_2 U3623 (.A1(data_i_10_), .A2(n4307), .B1(n3414), .Y(n3413));
sg13g2_nor2_2 U3624 (.A(n555), .B(n791), .Y(n3414));
sg13g2_inv_4 U3625 (.A(mixcol_data_o_10), .Y(n791));
sg13g2_inv_4 U3626 (.A(subbytes_data_o_10), .Y(n3409));
sg13g2_nor2_2 U3629 (.A(n3419), .B(n2248), .Y(n3418));
sg13g2_o21ai_1 U3630 (.A1(n4167), .A2(n3419), .B1(n3420), .Y(n3417));
sg13g2_nor2_2 U3632 (.A(n4165), .B(n793), .Y(n3422));
sg13g2_inv_4 U3633 (.A(n3421), .Y(n3415));
sg13g2_a21oi_2 U3635 (.A1(data_i_109_), .A2(n4307), .B1(n3424), .Y(n3423));
sg13g2_nor2_2 U3636 (.A(n555), .B(n793), .Y(n3424));
sg13g2_inv_4 U3637 (.A(mixcol_data_o_109), .Y(n793));
sg13g2_inv_4 U3638 (.A(subbytes_data_o_109), .Y(n3419));
sg13g2_o21ai_1 U3639 (.A1(n4332), .A2(n3425), .B1(n3426), .Y(addroundkey_data_i_108));
sg13g2_a21oi_2 U3640 (.A1(n4312), .A2(n3427), .B1(n3428), .Y(n3426));
sg13g2_nor2_2 U3641 (.A(n3429), .B(n2248), .Y(n3428));
sg13g2_o21ai_1 U3642 (.A1(n553), .A2(n3429), .B1(n3430), .Y(n3427));
sg13g2_a21oi_2 U3643 (.A1(n4315), .A2(n3431), .B1(n3432), .Y(n3430));
sg13g2_nor2_2 U3644 (.A(n4164), .B(n795), .Y(n3432));
sg13g2_inv_4 U3645 (.A(n3431), .Y(n3425));
sg13g2_o21ai_1 U3646 (.A1(n4327), .A2(n3429), .B1(n3433), .Y(n3431));
sg13g2_a21oi_2 U3647 (.A1(data_i_108_), .A2(n4307), .B1(n3434), .Y(n3433));
sg13g2_nor2_2 U3648 (.A(n555), .B(n795), .Y(n3434));
sg13g2_inv_4 U3649 (.A(mixcol_data_o_108), .Y(n795));
sg13g2_inv_4 U3650 (.A(subbytes_data_o_108), .Y(n3429));
sg13g2_o21ai_1 U3651 (.A1(n4332), .A2(n3435), .B1(n3436), .Y(addroundkey_data_i_107));
sg13g2_a21oi_2 U3652 (.A1(n4312), .A2(n3437), .B1(n3438), .Y(n3436));
sg13g2_nor2_2 U3653 (.A(n3439), .B(n2248), .Y(n3438));
sg13g2_o21ai_1 U3654 (.A1(n4167), .A2(n3439), .B1(n3440), .Y(n3437));
sg13g2_a21oi_2 U3655 (.A1(n4315), .A2(n3441), .B1(n3442), .Y(n3440));
sg13g2_nor2_2 U3656 (.A(n4164), .B(n797), .Y(n3442));
sg13g2_inv_4 U3657 (.A(n3441), .Y(n3435));
sg13g2_o21ai_1 U3658 (.A1(n4329), .A2(n3439), .B1(n3443), .Y(n3441));
sg13g2_a21oi_2 U3659 (.A1(data_i_107_), .A2(n4307), .B1(n3444), .Y(n3443));
sg13g2_nor2_2 U3660 (.A(n555), .B(n797), .Y(n3444));
sg13g2_inv_4 U3661 (.A(mixcol_data_o_107), .Y(n797));
sg13g2_inv_4 U3662 (.A(subbytes_data_o_107), .Y(n3439));
sg13g2_a21oi_2 U3664 (.A1(n4312), .A2(n3447), .B1(n3448), .Y(n3446));
sg13g2_nor2_2 U3665 (.A(n3449), .B(n2248), .Y(n3448));
sg13g2_o21ai_1 U3666 (.A1(n4167), .A2(n3449), .B1(n3450), .Y(n3447));
sg13g2_a21oi_2 U3667 (.A1(n4315), .A2(n3451), .B1(n3452), .Y(n3450));
sg13g2_nor2_2 U3668 (.A(n4165), .B(n799), .Y(n3452));
sg13g2_inv_4 U3669 (.A(n3451), .Y(n3445));
sg13g2_o21ai_1 U3670 (.A1(n4329), .A2(n3449), .B1(n3453), .Y(n3451));
sg13g2_a21oi_2 U3671 (.A1(data_i_106_), .A2(n4307), .B1(n3454), .Y(n3453));
sg13g2_nor2_2 U3672 (.A(n555), .B(n799), .Y(n3454));
sg13g2_inv_4 U3673 (.A(mixcol_data_o_106), .Y(n799));
sg13g2_inv_4 U3674 (.A(subbytes_data_o_106), .Y(n3449));
sg13g2_o21ai_1 U3675 (.A1(n4332), .A2(n3455), .B1(n3456), .Y(addroundkey_data_i_105));
sg13g2_a21oi_2 U3676 (.A1(n4312), .A2(n3457), .B1(n3458), .Y(n3456));
sg13g2_nor2_2 U3677 (.A(n3459), .B(n2248), .Y(n3458));
sg13g2_o21ai_1 U3678 (.A1(n553), .A2(n3459), .B1(n3460), .Y(n3457));
sg13g2_a21oi_2 U3679 (.A1(n4315), .A2(n3461), .B1(n3462), .Y(n3460));
sg13g2_nor2_2 U3680 (.A(n4165), .B(n801), .Y(n3462));
sg13g2_inv_4 U3681 (.A(n3461), .Y(n3455));
sg13g2_o21ai_1 U3682 (.A1(n4327), .A2(n3459), .B1(n3463), .Y(n3461));
sg13g2_a21oi_2 U3683 (.A1(data_i_105_), .A2(n4307), .B1(n3464), .Y(n3463));
sg13g2_nor2_2 U3684 (.A(n555), .B(n801), .Y(n3464));
sg13g2_inv_4 U3685 (.A(mixcol_data_o_105), .Y(n801));
sg13g2_inv_4 U3686 (.A(subbytes_data_o_105), .Y(n3459));
sg13g2_o21ai_1 U3687 (.A1(n4332), .A2(n3465), .B1(n3466), .Y(addroundkey_data_i_104));
sg13g2_a21oi_2 U3688 (.A1(n4312), .A2(n3467), .B1(n3468), .Y(n3466));
sg13g2_nor2_2 U3689 (.A(n3469), .B(n2248), .Y(n3468));
sg13g2_o21ai_1 U3690 (.A1(n4167), .A2(n3469), .B1(n3470), .Y(n3467));
sg13g2_a21oi_2 U3691 (.A1(n4315), .A2(n3471), .B1(n3472), .Y(n3470));
sg13g2_nor2_2 U3692 (.A(n4165), .B(n803), .Y(n3472));
sg13g2_inv_4 U3693 (.A(n3471), .Y(n3465));
sg13g2_o21ai_1 U3694 (.A1(n4330), .A2(n3469), .B1(n3473), .Y(n3471));
sg13g2_a21oi_2 U3695 (.A1(data_i_104_), .A2(n4307), .B1(n3474), .Y(n3473));
sg13g2_nor2_2 U3696 (.A(n555), .B(n803), .Y(n3474));
sg13g2_inv_4 U3697 (.A(mixcol_data_o_104), .Y(n803));
sg13g2_inv_4 U3698 (.A(subbytes_data_o_104), .Y(n3469));
sg13g2_o21ai_1 U3699 (.A1(n4332), .A2(n3475), .B1(n3476), .Y(addroundkey_data_i_103));
sg13g2_a21oi_2 U3700 (.A1(n4313), .A2(n3477), .B1(n3478), .Y(n3476));
sg13g2_nor2_2 U3701 (.A(n3479), .B(n2248), .Y(n3478));
sg13g2_o21ai_1 U3702 (.A1(n553), .A2(n3479), .B1(n3480), .Y(n3477));
sg13g2_a21oi_2 U3703 (.A1(n4315), .A2(n3481), .B1(n3482), .Y(n3480));
sg13g2_nor2_2 U3704 (.A(n4164), .B(n805), .Y(n3482));
sg13g2_inv_4 U3705 (.A(n3481), .Y(n3475));
sg13g2_o21ai_1 U3706 (.A1(n4328), .A2(n3479), .B1(n3483), .Y(n3481));
sg13g2_a21oi_2 U3707 (.A1(data_i_103_), .A2(n4307), .B1(n3484), .Y(n3483));
sg13g2_nor2_2 U3708 (.A(n555), .B(n805), .Y(n3484));
sg13g2_inv_4 U3709 (.A(mixcol_data_o_103), .Y(n805));
sg13g2_inv_4 U3710 (.A(subbytes_data_o_103), .Y(n3479));
sg13g2_o21ai_1 U3711 (.A1(n4332), .A2(n3485), .B1(n3486), .Y(addroundkey_data_i_102));
sg13g2_a21oi_2 U3712 (.A1(n4313), .A2(n3487), .B1(n3488), .Y(n3486));
sg13g2_nor2_2 U3713 (.A(n3489), .B(n2248), .Y(n3488));
sg13g2_o21ai_1 U3714 (.A1(n4167), .A2(n3489), .B1(n3490), .Y(n3487));
sg13g2_a21oi_2 U3715 (.A1(n4315), .A2(n3491), .B1(n3492), .Y(n3490));
sg13g2_nor2_2 U3716 (.A(n4164), .B(n807), .Y(n3492));
sg13g2_inv_4 U3717 (.A(n3491), .Y(n3485));
sg13g2_o21ai_1 U3718 (.A1(n4328), .A2(n3489), .B1(n3493), .Y(n3491));
sg13g2_a21oi_2 U3719 (.A1(data_i_102_), .A2(n4307), .B1(n3494), .Y(n3493));
sg13g2_nor2_2 U3720 (.A(n555), .B(n807), .Y(n3494));
sg13g2_inv_4 U3721 (.A(mixcol_data_o_102), .Y(n807));
sg13g2_inv_4 U3722 (.A(subbytes_data_o_102), .Y(n3489));
sg13g2_o21ai_1 U3723 (.A1(n4332), .A2(n3495), .B1(n3496), .Y(addroundkey_data_i_101));
sg13g2_a21oi_2 U3724 (.A1(n4313), .A2(n3497), .B1(n3498), .Y(n3496));
sg13g2_nor2_2 U3725 (.A(n3499), .B(n2248), .Y(n3498));
sg13g2_o21ai_1 U3726 (.A1(n4167), .A2(n3499), .B1(n3500), .Y(n3497));
sg13g2_a21oi_2 U3727 (.A1(n4315), .A2(n3501), .B1(n3502), .Y(n3500));
sg13g2_nor2_2 U3728 (.A(n4164), .B(n809), .Y(n3502));
sg13g2_inv_4 U3729 (.A(n3501), .Y(n3495));
sg13g2_o21ai_1 U3730 (.A1(n4330), .A2(n3499), .B1(n3503), .Y(n3501));
sg13g2_a21oi_2 U3731 (.A1(data_i_101_), .A2(n4307), .B1(n3504), .Y(n3503));
sg13g2_nor2_2 U3732 (.A(n555), .B(n809), .Y(n3504));
sg13g2_inv_4 U3733 (.A(mixcol_data_o_101), .Y(n809));
sg13g2_inv_4 U3734 (.A(subbytes_data_o_101), .Y(n3499));
sg13g2_o21ai_1 U3735 (.A1(n4332), .A2(n3505), .B1(n3506), .Y(addroundkey_data_i_100));
sg13g2_a21oi_2 U3736 (.A1(n4312), .A2(n3507), .B1(n3508), .Y(n3506));
sg13g2_nor2_2 U3737 (.A(n3509), .B(n2248), .Y(n3508));
sg13g2_o21ai_1 U3738 (.A1(n4167), .A2(n3509), .B1(n3510), .Y(n3507));
sg13g2_a21oi_2 U3739 (.A1(n4315), .A2(n3511), .B1(n3512), .Y(n3510));
sg13g2_nor2_2 U3740 (.A(n4164), .B(n811), .Y(n3512));
sg13g2_inv_4 U3741 (.A(n3511), .Y(n3505));
sg13g2_o21ai_1 U3742 (.A1(n4326), .A2(n3509), .B1(n3513), .Y(n3511));
sg13g2_a21oi_2 U3743 (.A1(data_i_100_), .A2(n4307), .B1(n3514), .Y(n3513));
sg13g2_nor2_2 U3744 (.A(n555), .B(n811), .Y(n3514));
sg13g2_inv_4 U3745 (.A(mixcol_data_o_100), .Y(n811));
sg13g2_inv_4 U3746 (.A(subbytes_data_o_100), .Y(n3509));
sg13g2_o21ai_1 U3747 (.A1(n4332), .A2(n3515), .B1(n3516), .Y(addroundkey_data_i_0));
sg13g2_a21oi_2 U3748 (.A1(n4313), .A2(n3517), .B1(n3518), .Y(n3516));
sg13g2_nor2_2 U3749 (.A(n3519), .B(n2248), .Y(n3518));
sg13g2_o21ai_1 U3751 (.A1(n553), .A2(n3519), .B1(n3521), .Y(n3517));
sg13g2_a21oi_2 U3752 (.A1(n4315), .A2(n3522), .B1(n3523), .Y(n3521));
sg13g2_nor2_2 U3753 (.A(n4165), .B(n813), .Y(n3523));
sg13g2_inv_4 U3760 (.A(n3522), .Y(n3515));
sg13g2_o21ai_1 U3761 (.A1(n4328), .A2(n3519), .B1(n3526), .Y(n3522));
sg13g2_a21oi_2 U3762 (.A1(data_i_0_), .A2(n4307), .B1(n3527), .Y(n3526));
sg13g2_nor2_2 U3763 (.A(n555), .B(n813), .Y(n3527));
sg13g2_inv_4 U3764 (.A(mixcol_data_o_0), .Y(n813));
sg13g2_inv_4 U3765 (.A(n1904), .Y(n2253));
sg13g2_inv_4 U3767 (.A(subbytes_data_o_0), .Y(n3519));
sg13g2_nand2_2 U3768 (.A(n4333), .B(n3528), .Y(N1567));
sg13g2_inv_4 U3769 (.A(n3529), .Y(N1566));
sg13g2_nor2_2 U3770 (.A(next_ready_o), .B(next_first_round_reg), .Y(n3529));
sg13g2_nor2_2 U3771 (.A(n3528), .B(n4332), .Y(next_first_round_reg));
sg13g2_inv_4 U3772 (.A(load_i), .Y(n3528));
sg13g2_nor2_2 U3773 (.A(n1118), .B(n4333), .Y(next_ready_o));
sg13g2_nand2_2 U3775 (.A(addroundkey_ready_o), .B(N587), .Y(n1118));
sg13g2_o21ai_1 U3779 (.A1(N1590), .A2(n3530), .B1(n3531), .Y(N1405));
sg13g2_nand2_2 U3780 (.A(N1590), .B(key_i_63_), .Y(n3531));
sg13g2_o21ai_1 U3782 (.A1(N1590), .A2(n3532), .B1(n3533), .Y(N1404));
sg13g2_nand2_2 U3783 (.A(N1590), .B(key_i_62_), .Y(n3533));
sg13g2_o21ai_1 U3785 (.A1(N1590), .A2(n3534), .B1(n3535), .Y(N1403));
sg13g2_nand2_2 U3786 (.A(N1590), .B(key_i_61_), .Y(n3535));
sg13g2_o21ai_1 U3788 (.A1(N1590), .A2(n3536), .B1(n3537), .Y(N1402));
sg13g2_nand2_2 U3789 (.A(N1590), .B(key_i_60_), .Y(n3537));
sg13g2_o21ai_1 U3791 (.A1(N1590), .A2(n3538), .B1(n3539), .Y(N1401));
sg13g2_nand2_2 U3792 (.A(N1590), .B(key_i_59_), .Y(n3539));
sg13g2_o21ai_1 U3794 (.A1(N1590), .A2(n3540), .B1(n3541), .Y(N1400));
sg13g2_nand2_2 U3795 (.A(N1590), .B(key_i_58_), .Y(n3541));
sg13g2_o21ai_1 U3797 (.A1(N1590), .A2(n3542), .B1(n3543), .Y(N1399));
sg13g2_nand2_2 U3798 (.A(N1590), .B(key_i_57_), .Y(n3543));
sg13g2_o21ai_1 U3800 (.A1(N1590), .A2(n3544), .B1(n3545), .Y(N1398));
sg13g2_nand2_2 U3801 (.A(N1590), .B(key_i_56_), .Y(n3545));
sg13g2_o21ai_1 U3803 (.A1(N1590), .A2(n3546), .B1(n3547), .Y(N1397));
sg13g2_nand2_2 U3804 (.A(N1590), .B(key_i_55_), .Y(n3547));
sg13g2_o21ai_1 U3806 (.A1(N1590), .A2(n3548), .B1(n3549), .Y(N1396));
sg13g2_nand2_2 U3807 (.A(N1590), .B(key_i_54_), .Y(n3549));
sg13g2_o21ai_1 U3809 (.A1(N1590), .A2(n3550), .B1(n3551), .Y(N1395));
sg13g2_nand2_2 U3810 (.A(N1590), .B(key_i_53_), .Y(n3551));
sg13g2_o21ai_1 U3812 (.A1(N1590), .A2(n3552), .B1(n3553), .Y(N1394));
sg13g2_nand2_2 U3813 (.A(N1590), .B(key_i_52_), .Y(n3553));
sg13g2_o21ai_1 U3815 (.A1(N1590), .A2(n3554), .B1(n3555), .Y(N1393));
sg13g2_nand2_2 U3816 (.A(N1590), .B(key_i_51_), .Y(n3555));
sg13g2_o21ai_1 U3818 (.A1(N1590), .A2(n3556), .B1(n3557), .Y(N1392));
sg13g2_nand2_2 U3819 (.A(N1590), .B(key_i_50_), .Y(n3557));
sg13g2_o21ai_1 U3821 (.A1(N1590), .A2(n3558), .B1(n3559), .Y(N1391));
sg13g2_nand2_2 U3822 (.A(N1590), .B(key_i_49_), .Y(n3559));
sg13g2_o21ai_1 U3824 (.A1(N1590), .A2(n3560), .B1(n3561), .Y(N1390));
sg13g2_nand2_2 U3825 (.A(N1590), .B(key_i_48_), .Y(n3561));
sg13g2_o21ai_1 U3827 (.A1(N1590), .A2(n3562), .B1(n3563), .Y(N1389));
sg13g2_nand2_2 U3828 (.A(N1590), .B(key_i_47_), .Y(n3563));
sg13g2_o21ai_1 U3830 (.A1(N1590), .A2(n3564), .B1(n3565), .Y(N1388));
sg13g2_nand2_2 U3831 (.A(N1590), .B(key_i_46_), .Y(n3565));
sg13g2_o21ai_1 U3833 (.A1(N1590), .A2(n3566), .B1(n3567), .Y(N1387));
sg13g2_nand2_2 U3834 (.A(N1590), .B(key_i_45_), .Y(n3567));
sg13g2_o21ai_1 U3836 (.A1(N1590), .A2(n3568), .B1(n3569), .Y(N1386));
sg13g2_nand2_2 U3837 (.A(N1590), .B(key_i_44_), .Y(n3569));
sg13g2_o21ai_1 U3839 (.A1(N1590), .A2(n3570), .B1(n3571), .Y(N1385));
sg13g2_nand2_2 U3840 (.A(N1590), .B(key_i_43_), .Y(n3571));
sg13g2_o21ai_1 U3842 (.A1(N1590), .A2(n3572), .B1(n3573), .Y(N1384));
sg13g2_nand2_2 U3843 (.A(N1590), .B(key_i_42_), .Y(n3573));
sg13g2_o21ai_1 U3845 (.A1(N1590), .A2(n3574), .B1(n3575), .Y(N1383));
sg13g2_nand2_2 U3846 (.A(N1590), .B(key_i_41_), .Y(n3575));
sg13g2_o21ai_1 U3848 (.A1(N1590), .A2(n3576), .B1(n3577), .Y(N1382));
sg13g2_nand2_2 U3849 (.A(N1590), .B(key_i_40_), .Y(n3577));
sg13g2_o21ai_1 U3851 (.A1(N1590), .A2(n3578), .B1(n3579), .Y(N1381));
sg13g2_nand2_2 U3852 (.A(N1590), .B(key_i_39_), .Y(n3579));
sg13g2_o21ai_1 U3854 (.A1(N1590), .A2(n3580), .B1(n3581), .Y(N1380));
sg13g2_nand2_2 U3855 (.A(N1590), .B(key_i_38_), .Y(n3581));
sg13g2_o21ai_1 U3857 (.A1(N1590), .A2(n3582), .B1(n3583), .Y(N1379));
sg13g2_nand2_2 U3858 (.A(N1590), .B(key_i_37_), .Y(n3583));
sg13g2_o21ai_1 U3860 (.A1(N1590), .A2(n3584), .B1(n3585), .Y(N1378));
sg13g2_nand2_2 U3861 (.A(N1590), .B(key_i_36_), .Y(n3585));
sg13g2_o21ai_1 U3863 (.A1(N1590), .A2(n3586), .B1(n3587), .Y(N1377));
sg13g2_nand2_2 U3864 (.A(N1590), .B(key_i_35_), .Y(n3587));
sg13g2_o21ai_1 U3866 (.A1(N1590), .A2(n3588), .B1(n3589), .Y(N1376));
sg13g2_nand2_2 U3867 (.A(N1590), .B(key_i_34_), .Y(n3589));
sg13g2_o21ai_1 U3869 (.A1(N1590), .A2(n3590), .B1(n3591), .Y(N1375));
sg13g2_nand2_2 U3870 (.A(N1590), .B(key_i_33_), .Y(n3591));
sg13g2_o21ai_1 U3872 (.A1(N1590), .A2(n3592), .B1(n3593), .Y(N1374));
sg13g2_nand2_2 U3873 (.A(N1590), .B(key_i_32_), .Y(n3593));
sg13g2_o21ai_1 U3875 (.A1(N1590), .A2(n3594), .B1(n3595), .Y(N1373));
sg13g2_nand2_2 U3876 (.A(N1590), .B(key_i_31_), .Y(n3595));
sg13g2_o21ai_1 U3878 (.A1(N1590), .A2(n3596), .B1(n3597), .Y(N1372));
sg13g2_nand2_2 U3879 (.A(N1590), .B(key_i_30_), .Y(n3597));
sg13g2_o21ai_1 U3881 (.A1(N1590), .A2(n3598), .B1(n3599), .Y(N1371));
sg13g2_nand2_2 U3882 (.A(N1590), .B(key_i_29_), .Y(n3599));
sg13g2_o21ai_1 U3884 (.A1(N1590), .A2(n3600), .B1(n3601), .Y(N1370));
sg13g2_nand2_2 U3885 (.A(N1590), .B(key_i_28_), .Y(n3601));
sg13g2_o21ai_1 U3887 (.A1(N1590), .A2(n3602), .B1(n3603), .Y(N1369));
sg13g2_nand2_2 U3888 (.A(N1590), .B(key_i_27_), .Y(n3603));
sg13g2_o21ai_1 U3890 (.A1(N1590), .A2(n3604), .B1(n3605), .Y(N1368));
sg13g2_nand2_2 U3891 (.A(N1590), .B(key_i_26_), .Y(n3605));
sg13g2_o21ai_1 U3893 (.A1(N1590), .A2(n3606), .B1(n3607), .Y(N1367));
sg13g2_nand2_2 U3894 (.A(N1590), .B(key_i_25_), .Y(n3607));
sg13g2_o21ai_1 U3896 (.A1(N1590), .A2(n3608), .B1(n3609), .Y(N1366));
sg13g2_nand2_2 U3897 (.A(N1590), .B(key_i_24_), .Y(n3609));
sg13g2_o21ai_1 U3899 (.A1(N1590), .A2(n3610), .B1(n3611), .Y(N1365));
sg13g2_nand2_2 U3900 (.A(N1590), .B(key_i_23_), .Y(n3611));
sg13g2_o21ai_1 U3902 (.A1(N1590), .A2(n3612), .B1(n3613), .Y(N1364));
sg13g2_nand2_2 U3903 (.A(N1590), .B(key_i_22_), .Y(n3613));
sg13g2_o21ai_1 U3905 (.A1(N1590), .A2(n3614), .B1(n3615), .Y(N1363));
sg13g2_nand2_2 U3906 (.A(N1590), .B(key_i_21_), .Y(n3615));
sg13g2_o21ai_1 U3908 (.A1(N1590), .A2(n3616), .B1(n3617), .Y(N1362));
sg13g2_nand2_2 U3909 (.A(N1590), .B(key_i_20_), .Y(n3617));
sg13g2_o21ai_1 U3911 (.A1(N1590), .A2(n3618), .B1(n3619), .Y(N1361));
sg13g2_nand2_2 U3912 (.A(N1590), .B(key_i_19_), .Y(n3619));
sg13g2_o21ai_1 U3914 (.A1(N1590), .A2(n3620), .B1(n3621), .Y(N1360));
sg13g2_nand2_2 U3915 (.A(N1590), .B(key_i_18_), .Y(n3621));
sg13g2_o21ai_1 U3917 (.A1(N1590), .A2(n3622), .B1(n3623), .Y(N1359));
sg13g2_nand2_2 U3918 (.A(N1590), .B(key_i_17_), .Y(n3623));
sg13g2_o21ai_1 U3920 (.A1(N1590), .A2(n3624), .B1(n3625), .Y(N1358));
sg13g2_nand2_2 U3921 (.A(N1590), .B(key_i_16_), .Y(n3625));
sg13g2_o21ai_1 U3923 (.A1(N1590), .A2(n3626), .B1(n3627), .Y(N1357));
sg13g2_nand2_2 U3924 (.A(N1590), .B(key_i_15_), .Y(n3627));
sg13g2_o21ai_1 U3926 (.A1(N1590), .A2(n3628), .B1(n3629), .Y(N1356));
sg13g2_nand2_2 U3927 (.A(N1590), .B(key_i_14_), .Y(n3629));
sg13g2_o21ai_1 U3929 (.A1(N1590), .A2(n3630), .B1(n3631), .Y(N1355));
sg13g2_nand2_2 U3930 (.A(N1590), .B(key_i_13_), .Y(n3631));
sg13g2_o21ai_1 U3932 (.A1(N1590), .A2(n3632), .B1(n3633), .Y(N1354));
sg13g2_nand2_2 U3933 (.A(N1590), .B(key_i_12_), .Y(n3633));
sg13g2_o21ai_1 U3935 (.A1(N1590), .A2(n3634), .B1(n3635), .Y(N1353));
sg13g2_nand2_2 U3936 (.A(N1590), .B(key_i_11_), .Y(n3635));
sg13g2_o21ai_1 U3938 (.A1(N1590), .A2(n3636), .B1(n3637), .Y(N1352));
sg13g2_nand2_2 U3939 (.A(N1590), .B(key_i_10_), .Y(n3637));
sg13g2_o21ai_1 U3941 (.A1(N1590), .A2(n3638), .B1(n3639), .Y(N1351));
sg13g2_nand2_2 U3942 (.A(N1590), .B(key_i_9_), .Y(n3639));
sg13g2_o21ai_1 U3944 (.A1(N1590), .A2(n3640), .B1(n3641), .Y(N1350));
sg13g2_nand2_2 U3945 (.A(N1590), .B(key_i_8_), .Y(n3641));
sg13g2_o21ai_1 U3947 (.A1(N1590), .A2(n3642), .B1(n3643), .Y(N1349));
sg13g2_nand2_2 U3948 (.A(N1590), .B(key_i_7_), .Y(n3643));
sg13g2_o21ai_1 U3950 (.A1(N1590), .A2(n3644), .B1(n3645), .Y(N1348));
sg13g2_nand2_2 U3951 (.A(N1590), .B(key_i_6_), .Y(n3645));
sg13g2_o21ai_1 U3953 (.A1(N1590), .A2(n3646), .B1(n3647), .Y(N1347));
sg13g2_nand2_2 U3954 (.A(N1590), .B(key_i_5_), .Y(n3647));
sg13g2_o21ai_1 U3956 (.A1(N1590), .A2(n3648), .B1(n3649), .Y(N1346));
sg13g2_nand2_2 U3957 (.A(N1590), .B(key_i_4_), .Y(n3649));
sg13g2_o21ai_1 U3959 (.A1(N1590), .A2(n3650), .B1(n3651), .Y(N1345));
sg13g2_nand2_2 U3960 (.A(N1590), .B(key_i_3_), .Y(n3651));
sg13g2_o21ai_1 U3962 (.A1(N1590), .A2(n3652), .B1(n3653), .Y(N1344));
sg13g2_nand2_2 U3963 (.A(N1590), .B(key_i_2_), .Y(n3653));
sg13g2_o21ai_1 U3965 (.A1(N1590), .A2(n3654), .B1(n3655), .Y(N1343));
sg13g2_nand2_2 U3966 (.A(N1590), .B(key_i_1_), .Y(n3655));
sg13g2_o21ai_1 U3968 (.A1(N1590), .A2(n3656), .B1(n3657), .Y(N1342));
sg13g2_nand2_2 U3969 (.A(N1590), .B(key_i_0_), .Y(n3657));
sg13g2_inv_4 U4004 (.A(n3691), .Y(N1625));
sg13g2_inv_4 U4007 (.A(n3694), .Y(N1628));
sg13g2_inv_4 U4008 (.A(n3695), .Y(N1125));
sg13g2_mux2_2 U4282 (.A0(addroundkey_round_3), .A1(next_addroundkey_round_3), .S(net24693), .X(n4136));
sg13g2_mux2_2 U4284 (.A0(last_key_half_63), .A1(next_last_key_half_63), .S(net24393), .X(n4135));
sg13g2_mux2_2 U4286 (.A0(data_o_127_), .A1(next_addroundkey_data_reg_127), .S(net24381), .X(n4134));
sg13g2_mux2_2 U4290 (.A0(n4332), .A1(n4333), .S(N1566), .X(n4132));
sg13g2_mux2_2 U4298 (.A0(data_o_0_), .A1(next_addroundkey_data_reg_0), .S(net24381), .X(n4128));
sg13g2_mux2_2 U4300 (.A0(data_o_1_), .A1(next_addroundkey_data_reg_1), .S(net24383), .X(n4127));
sg13g2_mux2_2 U4302 (.A0(data_o_2_), .A1(next_addroundkey_data_reg_2), .S(net24393), .X(n4126));
sg13g2_mux2_2 U4304 (.A0(data_o_3_), .A1(next_addroundkey_data_reg_3), .S(net24415), .X(n4125));
sg13g2_mux2_2 U4306 (.A0(data_o_4_), .A1(next_addroundkey_data_reg_4), .S(net24381), .X(n4124));
sg13g2_mux2_2 U4308 (.A0(data_o_5_), .A1(next_addroundkey_data_reg_5), .S(net24393), .X(n4123));
sg13g2_mux2_2 U4310 (.A0(data_o_6_), .A1(next_addroundkey_data_reg_6), .S(net24383), .X(n4122));
sg13g2_mux2_2 U4312 (.A0(data_o_7_), .A1(next_addroundkey_data_reg_7), .S(net24393), .X(n4121));
sg13g2_mux2_2 U4314 (.A0(data_o_8_), .A1(next_addroundkey_data_reg_8), .S(net24381), .X(n4120));
sg13g2_mux2_2 U4316 (.A0(data_o_9_), .A1(next_addroundkey_data_reg_9), .S(net24383), .X(n4119));
sg13g2_mux2_2 U4318 (.A0(data_o_10_), .A1(next_addroundkey_data_reg_10), .S(net24383), .X(n4118));
sg13g2_mux2_2 U4322 (.A0(data_o_12_), .A1(next_addroundkey_data_reg_12), .S(net24381), .X(n4116));
sg13g2_mux2_2 U4324 (.A0(data_o_13_), .A1(next_addroundkey_data_reg_13), .S(net24381), .X(n4115));
sg13g2_mux2_2 U4326 (.A0(data_o_14_), .A1(next_addroundkey_data_reg_14), .S(net24381), .X(n4114));
sg13g2_mux2_2 U4328 (.A0(data_o_15_), .A1(next_addroundkey_data_reg_15), .S(net24383), .X(n4113));
sg13g2_mux2_2 U4330 (.A0(data_o_16_), .A1(next_addroundkey_data_reg_16), .S(net24383), .X(n4112));
sg13g2_mux2_2 U4332 (.A0(data_o_17_), .A1(next_addroundkey_data_reg_17), .S(net24415), .X(n4111));
sg13g2_mux2_2 U4334 (.A0(data_o_18_), .A1(next_addroundkey_data_reg_18), .S(net24383), .X(n4110));
sg13g2_mux2_2 U4336 (.A0(data_o_19_), .A1(next_addroundkey_data_reg_19), .S(net24381), .X(n4109));
sg13g2_mux2_2 U4338 (.A0(data_o_20_), .A1(next_addroundkey_data_reg_20), .S(net24381), .X(n4108));
sg13g2_mux2_2 U4340 (.A0(data_o_21_), .A1(next_addroundkey_data_reg_21), .S(net24383), .X(n4107));
sg13g2_mux2_2 U4342 (.A0(data_o_22_), .A1(next_addroundkey_data_reg_22), .S(net24393), .X(n4106));
sg13g2_mux2_2 U4344 (.A0(data_o_23_), .A1(next_addroundkey_data_reg_23), .S(net24393), .X(n4105));
sg13g2_mux2_2 U4346 (.A0(data_o_24_), .A1(next_addroundkey_data_reg_24), .S(net24383), .X(n4104));
sg13g2_mux2_2 U4348 (.A0(data_o_25_), .A1(next_addroundkey_data_reg_25), .S(net24383), .X(n4103));
sg13g2_mux2_2 U4350 (.A0(data_o_26_), .A1(next_addroundkey_data_reg_26), .S(net24383), .X(n4102));
sg13g2_mux2_2 U4352 (.A0(data_o_27_), .A1(next_addroundkey_data_reg_27), .S(net24381), .X(n4101));
sg13g2_mux2_2 U4354 (.A0(data_o_28_), .A1(next_addroundkey_data_reg_28), .S(net24381), .X(n4100));
sg13g2_mux2_2 U4356 (.A0(data_o_29_), .A1(next_addroundkey_data_reg_29), .S(net24383), .X(n4099));
sg13g2_mux2_2 U4358 (.A0(data_o_30_), .A1(next_addroundkey_data_reg_30), .S(net24381), .X(n4098));
sg13g2_mux2_2 U4360 (.A0(data_o_31_), .A1(next_addroundkey_data_reg_31), .S(net24393), .X(n4097));
sg13g2_mux2_2 U4362 (.A0(data_o_32_), .A1(next_addroundkey_data_reg_32), .S(net24381), .X(n4096));
sg13g2_mux2_2 U4364 (.A0(data_o_33_), .A1(next_addroundkey_data_reg_33), .S(net24393), .X(n4095));
sg13g2_mux2_2 U4366 (.A0(data_o_34_), .A1(next_addroundkey_data_reg_34), .S(net24393), .X(n4094));
sg13g2_mux2_2 U4368 (.A0(data_o_35_), .A1(next_addroundkey_data_reg_35), .S(net24381), .X(n4093));
sg13g2_mux2_2 U4370 (.A0(data_o_36_), .A1(next_addroundkey_data_reg_36), .S(net24393), .X(n4092));
sg13g2_mux2_2 U4372 (.A0(data_o_37_), .A1(next_addroundkey_data_reg_37), .S(net24383), .X(n4091));
sg13g2_mux2_2 U4374 (.A0(data_o_38_), .A1(next_addroundkey_data_reg_38), .S(net24393), .X(n4090));
sg13g2_mux2_2 U4376 (.A0(data_o_39_), .A1(next_addroundkey_data_reg_39), .S(net24381), .X(n4089));
sg13g2_mux2_2 U4378 (.A0(data_o_40_), .A1(next_addroundkey_data_reg_40), .S(net24383), .X(n4088));
sg13g2_mux2_2 U4380 (.A0(data_o_41_), .A1(next_addroundkey_data_reg_41), .S(net24393), .X(n4087));
sg13g2_mux2_2 U4382 (.A0(data_o_42_), .A1(next_addroundkey_data_reg_42), .S(net24383), .X(n4086));
sg13g2_mux2_2 U4384 (.A0(data_o_43_), .A1(next_addroundkey_data_reg_43), .S(net24381), .X(n4085));
sg13g2_mux2_2 U4386 (.A0(data_o_44_), .A1(next_addroundkey_data_reg_44), .S(net24381), .X(n4084));
sg13g2_mux2_2 U4388 (.A0(data_o_45_), .A1(next_addroundkey_data_reg_45), .S(net24393), .X(n4083));
sg13g2_mux2_2 U4390 (.A0(data_o_46_), .A1(next_addroundkey_data_reg_46), .S(net24383), .X(n4082));
sg13g2_mux2_2 U4392 (.A0(data_o_47_), .A1(next_addroundkey_data_reg_47), .S(net24381), .X(n4081));
sg13g2_mux2_2 U4394 (.A0(data_o_48_), .A1(next_addroundkey_data_reg_48), .S(net24393), .X(n4080));
sg13g2_mux2_2 U4396 (.A0(data_o_49_), .A1(next_addroundkey_data_reg_49), .S(net24393), .X(n4079));
sg13g2_mux2_2 U4398 (.A0(data_o_50_), .A1(next_addroundkey_data_reg_50), .S(net24393), .X(n4078));
sg13g2_mux2_2 U4400 (.A0(data_o_51_), .A1(next_addroundkey_data_reg_51), .S(net24381), .X(n4077));
sg13g2_mux2_2 U4402 (.A0(data_o_52_), .A1(next_addroundkey_data_reg_52), .S(net24381), .X(n4076));
sg13g2_mux2_2 U4404 (.A0(data_o_53_), .A1(next_addroundkey_data_reg_53), .S(net24393), .X(n4075));
sg13g2_mux2_2 U4406 (.A0(data_o_54_), .A1(next_addroundkey_data_reg_54), .S(net24383), .X(n4074));
sg13g2_mux2_2 U4408 (.A0(data_o_55_), .A1(next_addroundkey_data_reg_55), .S(net24383), .X(n4073));
sg13g2_mux2_2 U4410 (.A0(data_o_56_), .A1(next_addroundkey_data_reg_56), .S(net24393), .X(n4072));
sg13g2_mux2_2 U4412 (.A0(data_o_57_), .A1(next_addroundkey_data_reg_57), .S(net24393), .X(n4071));
sg13g2_mux2_2 U4414 (.A0(data_o_58_), .A1(next_addroundkey_data_reg_58), .S(net24393), .X(n4070));
sg13g2_mux2_2 U4416 (.A0(data_o_59_), .A1(next_addroundkey_data_reg_59), .S(net24393), .X(n4069));
sg13g2_mux2_2 U4418 (.A0(data_o_60_), .A1(next_addroundkey_data_reg_60), .S(net24393), .X(n4068));
sg13g2_mux2_2 U4420 (.A0(data_o_61_), .A1(next_addroundkey_data_reg_61), .S(net24393), .X(n4067));
sg13g2_mux2_2 U4422 (.A0(data_o_62_), .A1(next_addroundkey_data_reg_62), .S(net24393), .X(n4066));
sg13g2_mux2_2 U4424 (.A0(data_o_63_), .A1(next_addroundkey_data_reg_63), .S(net24393), .X(n4065));
sg13g2_mux2_2 U4426 (.A0(data_o_64_), .A1(next_addroundkey_data_reg_64), .S(net24393), .X(n4064));
sg13g2_mux2_2 U4428 (.A0(data_o_65_), .A1(next_addroundkey_data_reg_65), .S(net24393), .X(n4063));
sg13g2_mux2_2 U4430 (.A0(data_o_66_), .A1(next_addroundkey_data_reg_66), .S(net24393), .X(n4062));
sg13g2_mux2_2 U4432 (.A0(data_o_67_), .A1(next_addroundkey_data_reg_67), .S(net24393), .X(n4061));
sg13g2_mux2_2 U4434 (.A0(data_o_68_), .A1(next_addroundkey_data_reg_68), .S(net24393), .X(n4060));
sg13g2_mux2_2 U4436 (.A0(data_o_69_), .A1(next_addroundkey_data_reg_69), .S(net24393), .X(n4059));
sg13g2_mux2_2 U4438 (.A0(data_o_70_), .A1(next_addroundkey_data_reg_70), .S(net24383), .X(n4058));
sg13g2_mux2_2 U4440 (.A0(data_o_71_), .A1(next_addroundkey_data_reg_71), .S(net24415), .X(n4057));
sg13g2_mux2_2 U4442 (.A0(data_o_72_), .A1(next_addroundkey_data_reg_72), .S(net24381), .X(n4056));
sg13g2_mux2_2 U4446 (.A0(data_o_74_), .A1(next_addroundkey_data_reg_74), .S(net24381), .X(n4054));
sg13g2_mux2_2 U4448 (.A0(data_o_75_), .A1(next_addroundkey_data_reg_75), .S(net24415), .X(n4053));
sg13g2_mux2_2 U4450 (.A0(data_o_76_), .A1(next_addroundkey_data_reg_76), .S(net24383), .X(n4052));
sg13g2_mux2_2 U4452 (.A0(data_o_77_), .A1(next_addroundkey_data_reg_77), .S(net24415), .X(n4051));
sg13g2_mux2_2 U4454 (.A0(data_o_78_), .A1(next_addroundkey_data_reg_78), .S(net24383), .X(n4050));
sg13g2_mux2_2 U4456 (.A0(data_o_79_), .A1(next_addroundkey_data_reg_79), .S(net24383), .X(n4049));
sg13g2_mux2_2 U4458 (.A0(data_o_80_), .A1(next_addroundkey_data_reg_80), .S(net24393), .X(n4048));
sg13g2_mux2_2 U4460 (.A0(data_o_81_), .A1(next_addroundkey_data_reg_81), .S(net24381), .X(n4047));
sg13g2_mux2_2 U4462 (.A0(data_o_82_), .A1(next_addroundkey_data_reg_82), .S(net24383), .X(n4046));
sg13g2_mux2_2 U4464 (.A0(data_o_83_), .A1(next_addroundkey_data_reg_83), .S(net24383), .X(n4045));
sg13g2_mux2_2 U4466 (.A0(data_o_84_), .A1(next_addroundkey_data_reg_84), .S(net24383), .X(n4044));
sg13g2_mux2_2 U4468 (.A0(data_o_85_), .A1(next_addroundkey_data_reg_85), .S(net24393), .X(n4043));
sg13g2_mux2_2 U4470 (.A0(data_o_86_), .A1(next_addroundkey_data_reg_86), .S(net24381), .X(n4042));
sg13g2_mux2_2 U4472 (.A0(data_o_87_), .A1(next_addroundkey_data_reg_87), .S(net24415), .X(n4041));
sg13g2_mux2_2 U4474 (.A0(data_o_88_), .A1(next_addroundkey_data_reg_88), .S(net24393), .X(n4040));
sg13g2_mux2_2 U4476 (.A0(data_o_89_), .A1(next_addroundkey_data_reg_89), .S(net24381), .X(n4039));
sg13g2_mux2_2 U4478 (.A0(data_o_90_), .A1(next_addroundkey_data_reg_90), .S(net24381), .X(n4038));
sg13g2_mux2_2 U4480 (.A0(data_o_91_), .A1(next_addroundkey_data_reg_91), .S(net24393), .X(n4037));
sg13g2_mux2_2 U4482 (.A0(data_o_92_), .A1(next_addroundkey_data_reg_92), .S(net24393), .X(n4036));
sg13g2_mux2_2 U4484 (.A0(data_o_93_), .A1(next_addroundkey_data_reg_93), .S(net24393), .X(n4035));
sg13g2_mux2_2 U4486 (.A0(data_o_94_), .A1(next_addroundkey_data_reg_94), .S(net24393), .X(n4034));
sg13g2_mux2_2 U4488 (.A0(data_o_95_), .A1(next_addroundkey_data_reg_95), .S(net24383), .X(n4033));
sg13g2_mux2_2 U4490 (.A0(data_o_96_), .A1(next_addroundkey_data_reg_96), .S(net24383), .X(n4032));
sg13g2_mux2_2 U4492 (.A0(data_o_97_), .A1(next_addroundkey_data_reg_97), .S(net24383), .X(n4031));
sg13g2_mux2_2 U4494 (.A0(data_o_98_), .A1(next_addroundkey_data_reg_98), .S(net24383), .X(n4030));
sg13g2_mux2_2 U4498 (.A0(data_o_99_), .A1(next_addroundkey_data_reg_99), .S(net24381), .X(n4028));
sg13g2_mux2_2 U4500 (.A0(data_o_100_), .A1(next_addroundkey_data_reg_100), .S(net24393), .X(n4027));
sg13g2_mux2_2 U4502 (.A0(data_o_101_), .A1(next_addroundkey_data_reg_101), .S(net24415), .X(n4026));
sg13g2_mux2_2 U4504 (.A0(data_o_102_), .A1(next_addroundkey_data_reg_102), .S(net24381), .X(n4025));
sg13g2_mux2_2 U4506 (.A0(data_o_103_), .A1(next_addroundkey_data_reg_103), .S(net24381), .X(n4024));
sg13g2_mux2_2 U4508 (.A0(data_o_104_), .A1(next_addroundkey_data_reg_104), .S(net24383), .X(n4023));
sg13g2_mux2_2 U4510 (.A0(data_o_105_), .A1(next_addroundkey_data_reg_105), .S(net24383), .X(n4022));
sg13g2_mux2_2 U4512 (.A0(data_o_106_), .A1(next_addroundkey_data_reg_106), .S(net24381), .X(n4021));
sg13g2_mux2_2 U4514 (.A0(data_o_107_), .A1(next_addroundkey_data_reg_107), .S(net24381), .X(n4020));
sg13g2_mux2_2 U4516 (.A0(data_o_108_), .A1(next_addroundkey_data_reg_108), .S(net24383), .X(n4019));
sg13g2_mux2_2 U4518 (.A0(data_o_109_), .A1(next_addroundkey_data_reg_109), .S(net24381), .X(n4018));
sg13g2_mux2_2 U4520 (.A0(data_o_110_), .A1(next_addroundkey_data_reg_110), .S(net24393), .X(n4017));
sg13g2_mux2_2 U4522 (.A0(data_o_111_), .A1(next_addroundkey_data_reg_111), .S(net24381), .X(n4016));
sg13g2_mux2_2 U4524 (.A0(data_o_112_), .A1(next_addroundkey_data_reg_112), .S(net24381), .X(n4015));
sg13g2_mux2_2 U4526 (.A0(data_o_113_), .A1(next_addroundkey_data_reg_113), .S(net24383), .X(n4014));
sg13g2_mux2_2 U4528 (.A0(data_o_114_), .A1(next_addroundkey_data_reg_114), .S(net24393), .X(n4013));
sg13g2_mux2_2 U4530 (.A0(data_o_115_), .A1(next_addroundkey_data_reg_115), .S(net24383), .X(n4012));
sg13g2_mux2_2 U4532 (.A0(data_o_116_), .A1(next_addroundkey_data_reg_116), .S(net24383), .X(n4011));
sg13g2_mux2_2 U4534 (.A0(data_o_117_), .A1(next_addroundkey_data_reg_117), .S(net24383), .X(n4010));
sg13g2_mux2_2 U4536 (.A0(data_o_118_), .A1(next_addroundkey_data_reg_118), .S(net24383), .X(n4009));
sg13g2_mux2_2 U4538 (.A0(data_o_119_), .A1(next_addroundkey_data_reg_119), .S(net24383), .X(n4008));
sg13g2_mux2_2 U4540 (.A0(data_o_120_), .A1(next_addroundkey_data_reg_120), .S(net24383), .X(n4007));
sg13g2_mux2_2 U4542 (.A0(data_o_121_), .A1(next_addroundkey_data_reg_121), .S(net24383), .X(n4006));
sg13g2_mux2_2 U4544 (.A0(data_o_122_), .A1(next_addroundkey_data_reg_122), .S(net24383), .X(n4005));
sg13g2_mux2_2 U4546 (.A0(data_o_123_), .A1(next_addroundkey_data_reg_123), .S(net24383), .X(n4004));
sg13g2_mux2_2 U4548 (.A0(data_o_124_), .A1(next_addroundkey_data_reg_124), .S(net24383), .X(n4003));
sg13g2_mux2_2 U4550 (.A0(data_o_125_), .A1(next_addroundkey_data_reg_125), .S(net24383), .X(n4002));
sg13g2_mux2_2 U4552 (.A0(data_o_126_), .A1(next_addroundkey_data_reg_126), .S(net24383), .X(n4001));
sg13g2_mux2_2 U4554 (.A0(last_key_half_0), .A1(next_last_key_half_0), .S(net24383), .X(n4000));
sg13g2_mux2_2 U4556 (.A0(last_key_half_1), .A1(next_last_key_half_1), .S(net24383), .X(n3999));
sg13g2_mux2_2 U4558 (.A0(last_key_half_2), .A1(next_last_key_half_2), .S(net24381), .X(n3998));
sg13g2_mux2_2 U4560 (.A0(last_key_half_3), .A1(next_last_key_half_3), .S(net24381), .X(n3997));
sg13g2_mux2_2 U4562 (.A0(last_key_half_4), .A1(next_last_key_half_4), .S(net24381), .X(n3996));
sg13g2_mux2_2 U4564 (.A0(last_key_half_5), .A1(next_last_key_half_5), .S(net24381), .X(n3995));
sg13g2_mux2_2 U4566 (.A0(last_key_half_6), .A1(next_last_key_half_6), .S(net24381), .X(n3994));
sg13g2_mux2_2 U4568 (.A0(last_key_half_7), .A1(next_last_key_half_7), .S(net24381), .X(n3993));
sg13g2_mux2_2 U4570 (.A0(last_key_half_8), .A1(next_last_key_half_8), .S(net24381), .X(n3992));
sg13g2_mux2_2 U4572 (.A0(last_key_half_9), .A1(next_last_key_half_9), .S(net24381), .X(n3991));
sg13g2_mux2_2 U4574 (.A0(last_key_half_10), .A1(next_last_key_half_10), .S(net24381), .X(n3990));
sg13g2_mux2_2 U4576 (.A0(last_key_half_11), .A1(next_last_key_half_11), .S(net24381), .X(n3989));
sg13g2_mux2_2 U4578 (.A0(last_key_half_12), .A1(next_last_key_half_12), .S(net24381), .X(n3988));
sg13g2_mux2_2 U4580 (.A0(last_key_half_13), .A1(next_last_key_half_13), .S(net24381), .X(n3987));
sg13g2_mux2_2 U4582 (.A0(last_key_half_14), .A1(next_last_key_half_14), .S(net24381), .X(n3986));
sg13g2_mux2_2 U4584 (.A0(last_key_half_15), .A1(next_last_key_half_15), .S(net24381), .X(n3985));
sg13g2_mux2_2 U4586 (.A0(last_key_half_16), .A1(next_last_key_half_16), .S(net24383), .X(n3984));
sg13g2_mux2_2 U4588 (.A0(last_key_half_17), .A1(next_last_key_half_17), .S(net24383), .X(n3983));
sg13g2_mux2_2 U4590 (.A0(last_key_half_18), .A1(next_last_key_half_18), .S(net24381), .X(n3982));
sg13g2_mux2_2 U4592 (.A0(last_key_half_19), .A1(next_last_key_half_19), .S(net24381), .X(n3981));
sg13g2_mux2_2 U4594 (.A0(last_key_half_20), .A1(next_last_key_half_20), .S(net24383), .X(n3980));
sg13g2_mux2_2 U4596 (.A0(last_key_half_21), .A1(next_last_key_half_21), .S(net24383), .X(n3979));
sg13g2_mux2_2 U4598 (.A0(last_key_half_22), .A1(next_last_key_half_22), .S(net24381), .X(n3978));
sg13g2_mux2_2 U4600 (.A0(last_key_half_23), .A1(next_last_key_half_23), .S(net24393), .X(n3977));
sg13g2_mux2_2 U4602 (.A0(last_key_half_24), .A1(next_last_key_half_24), .S(net24383), .X(n3976));
sg13g2_mux2_2 U4604 (.A0(last_key_half_25), .A1(next_last_key_half_25), .S(net24381), .X(n3975));
sg13g2_mux2_2 U4606 (.A0(last_key_half_26), .A1(next_last_key_half_26), .S(net24383), .X(n3974));
sg13g2_mux2_2 U4608 (.A0(last_key_half_27), .A1(next_last_key_half_27), .S(net24393), .X(n3973));
sg13g2_mux2_2 U4612 (.A0(last_key_half_29), .A1(next_last_key_half_29), .S(net24383), .X(n3971));
sg13g2_mux2_2 U4614 (.A0(last_key_half_30), .A1(next_last_key_half_30), .S(net24393), .X(n3970));
sg13g2_mux2_2 U4616 (.A0(last_key_half_31), .A1(next_last_key_half_31), .S(net24381), .X(n3969));
sg13g2_mux2_2 U4618 (.A0(last_key_half_32), .A1(next_last_key_half_32), .S(net24381), .X(n3968));
sg13g2_mux2_2 U4620 (.A0(last_key_half_33), .A1(next_last_key_half_33), .S(net24393), .X(n3967));
sg13g2_mux2_2 U4622 (.A0(last_key_half_34), .A1(next_last_key_half_34), .S(net24383), .X(n3966));
sg13g2_mux2_2 U4624 (.A0(last_key_half_35), .A1(next_last_key_half_35), .S(net24383), .X(n3965));
sg13g2_mux2_2 U4626 (.A0(last_key_half_36), .A1(next_last_key_half_36), .S(net24393), .X(n3964));
sg13g2_mux2_2 U4628 (.A0(last_key_half_37), .A1(next_last_key_half_37), .S(net24381), .X(n3963));
sg13g2_mux2_2 U4630 (.A0(last_key_half_38), .A1(next_last_key_half_38), .S(net24393), .X(n3962));
sg13g2_mux2_2 U4632 (.A0(last_key_half_39), .A1(next_last_key_half_39), .S(net24383), .X(n3961));
sg13g2_mux2_2 U4634 (.A0(last_key_half_40), .A1(next_last_key_half_40), .S(net24381), .X(n3960));
sg13g2_mux2_2 U4636 (.A0(last_key_half_41), .A1(next_last_key_half_41), .S(net24393), .X(n3959));
sg13g2_mux2_2 U4638 (.A0(last_key_half_42), .A1(next_last_key_half_42), .S(net24393), .X(n3958));
sg13g2_mux2_2 U4640 (.A0(last_key_half_43), .A1(next_last_key_half_43), .S(net24381), .X(n3957));
sg13g2_mux2_2 U4642 (.A0(last_key_half_44), .A1(next_last_key_half_44), .S(net24393), .X(n3956));
sg13g2_mux2_2 U4644 (.A0(last_key_half_45), .A1(next_last_key_half_45), .S(net24383), .X(n3955));
sg13g2_mux2_2 U4646 (.A0(last_key_half_46), .A1(next_last_key_half_46), .S(net24393), .X(n3954));
sg13g2_mux2_2 U4648 (.A0(last_key_half_47), .A1(next_last_key_half_47), .S(net24393), .X(n3953));
sg13g2_mux2_2 U4650 (.A0(last_key_half_48), .A1(next_last_key_half_48), .S(net24381), .X(n3952));
sg13g2_mux2_2 U4654 (.A0(last_key_half_50), .A1(next_last_key_half_50), .S(net24383), .X(n3950));
sg13g2_mux2_2 U4656 (.A0(last_key_half_51), .A1(next_last_key_half_51), .S(net24393), .X(n3949));
sg13g2_mux2_2 U4658 (.A0(last_key_half_52), .A1(next_last_key_half_52), .S(net24393), .X(n3948));
sg13g2_mux2_2 U4660 (.A0(last_key_half_53), .A1(next_last_key_half_53), .S(net24381), .X(n3947));
sg13g2_mux2_2 U4662 (.A0(last_key_half_54), .A1(next_last_key_half_54), .S(net24381), .X(n3946));
sg13g2_mux2_2 U4664 (.A0(last_key_half_55), .A1(next_last_key_half_55), .S(net24381), .X(n3945));
sg13g2_mux2_2 U4666 (.A0(last_key_half_56), .A1(next_last_key_half_56), .S(net24383), .X(n3944));
sg13g2_mux2_2 U4668 (.A0(last_key_half_57), .A1(next_last_key_half_57), .S(net24381), .X(n3943));
sg13g2_mux2_2 U4670 (.A0(last_key_half_58), .A1(next_last_key_half_58), .S(net24393), .X(n3942));
sg13g2_mux2_2 U4672 (.A0(last_key_half_59), .A1(next_last_key_half_59), .S(net24383), .X(n3941));
sg13g2_mux2_2 U4674 (.A0(last_key_half_60), .A1(next_last_key_half_60), .S(net24393), .X(n3940));
sg13g2_mux2_2 U4676 (.A0(last_key_half_61), .A1(next_last_key_half_61), .S(net24383), .X(n3939));
sg13g2_mux2_2 U4678 (.A0(addroundkey_round_0), .A1(next_addroundkey_round_0), .S(net24693), .X(n3938));
sg13g2_mux2_2 U4680 (.A0(addroundkey_round_1), .A1(next_addroundkey_round_1), .S(net24693), .X(n3937));
sg13g2_mux2_2 U4682 (.A0(addroundkey_round_2), .A1(next_addroundkey_round_2), .S(net24693), .X(n3936));
sg13g2_nand2_2 U4686 (.A(r371_n27), .B(net25972), .Y(n4137));
sg13g2_xnor2_1 U4687 (.A(n4137), .B(net26538), .Y(N174));
sg13g2_inv_4 U4688 (.A(n4137), .Y(n4138));
sg13g2_nand2_2 U4689 (.A(net26538), .B(n4138), .Y(n4139));
sg13g2_xnor2_1 U4690 (.A(n4139), .B(net47654), .Y(N175));
sg13g2_nand2_2 U4718 (.A(addroundkey_round_1), .B(addroundkey_round_0), .Y(n4152));
sg13g2_xnor2_1 U4719 (.A(n4152), .B(addroundkey_round_2), .Y(N1537));
sg13g2_inv_4 U4720 (.A(n4152), .Y(n4153));
sg13g2_nand2_2 U4721 (.A(addroundkey_round_2), .B(n4153), .Y(n4154));
sg13g2_xnor2_1 U4722 (.A(n4154), .B(addroundkey_round_3), .Y(N1538));
sg13g2_o21ai_1 U4723 (.A1(net24787), .A2(n1042), .B1(n2035), .Y(keysched_last_key_i_24));
sg13g2_o21ai_1 U4724 (.A1(n1026), .A2(net24787), .B1(n2031), .Y(keysched_last_key_i_28));
sg13g2_inv_4 U4725 (.A(net24821), .Y(net24801));
sg13g2_o21ai_1 U4726 (.A1(net24783), .A2(n1090), .B1(n2151), .Y(keysched_last_key_i_13));
sg13g2_nand2_2 U4727 (.A(n4216), .B(n2235), .Y(keysched_last_key_i_0));
sg13g2_inv_4 U4728 (.A(net25885), .Y(net26430));
sg13g2_buf_8 U4729 (.A(net24863), .X(n4155));
sg13g2_nand2_2 U4730 (.A(n4233), .B(key_i_11_), .Y(n4270));
sg13g2_inv_4 U4731 (.A(net24823), .Y(net24791));
sg13g2_nand2_2 U4732 (.A(n4215), .B(key_i_0_), .Y(n4216));
sg13g2_nand2_2 U4733 (.A(net24821), .B(key_i_1_), .Y(n4299));
sg13g2_inv_4 U4734 (.A(net25885), .Y(n4156));
sg13g2_inv_4 U4735 (.A(net25885), .Y(n4239));
sg13g2_inv_4 U4736 (.A(net26049), .Y(net24839));
sg13g2_inv_4 U4737 (.A(net24881), .Y(net26049));
sg13g2_nand2_2 U4738 (.A(keysched_new_key_o_9), .B(net24839), .Y(n4235));
sg13g2_inv_4 U4739 (.A(net26210), .Y(n4233));
sg13g2_nand2_2 U4740 (.A(net24879), .B(keysched_new_key_o_4), .Y(n2007));
sg13g2_nand2_2 U4741 (.A(n168), .B(n4158), .Y(n4159));
sg13g2_inv_4 U4742 (.A(net26078), .Y(n4157));
sg13g2_inv_4 U4743 (.A(n4277), .Y(n4158));
sg13g2_inv_4 U4744 (.A(n4159), .Y(n4160));
sg13g2_nand2_2 U4745 (.A(n4157), .B(n4158), .Y(n4161));
sg13g2_nand3_1 U4746 (.A(net27301), .B(n4210), .C(n4228), .Y(net26078));
sg13g2_inv_4 U4747 (.A(net24825), .Y(net24821));
sg13g2_o21ai_1 U4748 (.A1(net26188), .A2(n2175), .B1(n2176), .Y(keysched_last_key_i_128));
sg13g2_inv_4 U4749 (.A(net24633), .Y(net24611));
sg13g2_inv_4 U4750 (.A(n4282), .Y(net24633));
sg13g2_nand2_2 U4751 (.A(N1613), .B(decrypt_i), .Y(n4162));
sg13g2_inv_4 U4752 (.A(n2248), .Y(n4311));
sg13g2_inv_4 U4753 (.A(n560), .Y(n4163));
sg13g2_inv_4 U4754 (.A(sbox_data_o_7), .Y(n4268));
sg13g2_inv_4 U4755 (.A(n4163), .Y(n4323));
sg13g2_o21ai_1 U4756 (.A1(n4221), .A2(n2099), .B1(n2100), .Y(keysched_last_key_i_164));
sg13g2_inv_4 U4757 (.A(n4296), .Y(n555));
sg13g2_inv_4 U4758 (.A(n4284), .Y(n4296));
sg13g2_a21oi_2 U4759 (.A1(n2244), .A2(n2917), .B1(n2918), .Y(n2916));
sg13g2_nand4_1 U4760 (.A(n4161), .B(n4282), .C(n4283), .D(n4281), .Y(n857));
sg13g2_mux2_2 U4761 (.A0(last_key_half_49), .A1(next_last_key_half_49), .S(net24393), .X(n3951));
sg13g2_inv_4 U4762 (.A(n1912), .Y(net27141));
sg13g2_nand2_2 U4763 (.A(N29), .B(mixcol_ready_o), .Y(n4164));
sg13g2_nand2_2 U4764 (.A(N29), .B(mixcol_ready_o), .Y(n4165));
sg13g2_o21ai_1 U4765 (.A1(n4221), .A2(n2097), .B1(n2098), .Y(keysched_last_key_i_165));
sg13g2_inv_4 U4766 (.A(sbox_data_o_2), .Y(n4226));
sg13g2_inv_4 U4767 (.A(net24823), .Y(net24795));
sg13g2_inv_4 U4768 (.A(net26302), .Y(net24823));
sg13g2_inv_4 U4769 (.A(n4215), .Y(n4211));
sg13g2_nand2_2 U4770 (.A(decrypt_i), .B(subbytes_ready_o), .Y(n4166));
sg13g2_nand2_2 U4771 (.A(decrypt_i), .B(subbytes_ready_o), .Y(n4167));
sg13g2_nand2_2 U4772 (.A(decrypt_i), .B(subbytes_ready_o), .Y(n553));
sg13g2_o21ai_1 U4773 (.A1(net26188), .A2(n2110), .B1(n2111), .Y(keysched_last_key_i_159));
sg13g2_o21ai_1 U4774 (.A1(n4221), .A2(n2059), .B1(n2060), .Y(keysched_last_key_i_183));
sg13g2_o21ai_1 U4775 (.A1(net24801), .A2(n2105), .B1(n2106), .Y(keysched_last_key_i_161));
sg13g2_o21ai_1 U4776 (.A1(n974), .A2(net24825), .B1(n2018), .Y(keysched_last_key_i_3));
sg13g2_nand2_2 U4777 (.A(N1659), .B(keysched_ready_o), .Y(net39126));
sg13g2_nand2_2 U4778 (.A(net44478), .B(n4174), .Y(n4170));
sg13g2_nand2_2 U4779 (.A(n4170), .B(n4171), .Y(n4168));
sg13g2_inv_4 U4780 (.A(n4168), .Y(n4256));
sg13g2_nor2_2 U4781 (.A(n4172), .B(net44473), .Y(n4169));
sg13g2_inv_4 U4782 (.A(n4169), .Y(n4171));
sg13g2_inv_4 U4783 (.A(N1559), .Y(n4172));
sg13g2_nand2_2 U4784 (.A(net43702), .B(N1559), .Y(n4173));
sg13g2_inv_4 U4785 (.A(n4173), .Y(n4174));
sg13g2_inv_4 U4786 (.A(net24827), .Y(n4215));
sg13g2_nand3_1 U4787 (.A(net27301), .B(n4210), .C(n4228), .Y(n4175));
sg13g2_xnor2_1 U4788 (.A(three_2), .B(net44332), .Y(r372_n15));
sg13g2_nand2_2 U4789 (.A(N1645), .B(keysched_ready_o), .Y(n4219));
sg13g2_o21ai_1 U4790 (.A1(n4328), .A2(n595), .B1(n596), .Y(subbytes_data_i_83));
sg13g2_xnor2_1 U4791 (.A(net47651), .B(net26537), .Y(four_3_));
sg13g2_xnor2_1 U4792 (.A(N7), .B(addroundkey_round_1), .Y(r373_n17));
sg13g2_inv_4 U4793 (.A(n1131), .Y(net26981));
sg13g2_inv_4 U4794 (.A(n4212), .Y(n4213));
sg13g2_o21ai_1 U4795 (.A1(n4221), .A2(n2063), .B1(n2064), .Y(keysched_last_key_i_181));
sg13g2_a21oi_2 U4796 (.A1(state), .A2(N587), .B1(n557), .Y(subbytes_start_i));
sg13g2_o21ai_1 U4797 (.A1(net24693), .A2(n946), .B1(n947), .Y(next_last_key_half_46));
sg13g2_nand2_2 U4798 (.A(n4323), .B(data_o_78_), .Y(n608));
sg13g2_nor2_2 U4799 (.A(n4176), .B(net44654), .Y(net44818));
sg13g2_inv_4 U4800 (.A(net26019), .Y(n4176));
sg13g2_nand2_2 U4801 (.A(n4323), .B(data_o_86_), .Y(n590));
sg13g2_nand2_2 U4802 (.A(addroundkey_round_3), .B(n4272), .Y(n4271));
sg13g2_nand2_2 U4803 (.A(n4323), .B(data_o_118_), .Y(n774));
sg13g2_nand4_1 U4804 (.A(net26537), .B(N7), .C(three_0), .D(net47651), .Y(N1610));
sg13g2_inv_4 U4805 (.A(net25928), .Y(N7));
sg13g2_o21ai_1 U4806 (.A1(net44819), .A2(n4177), .B1(net44320), .Y(n4272));
sg13g2_inv_4 U4807 (.A(n168), .Y(n4177));
sg13g2_nand2_2 U4808 (.A(n3525), .B(n843), .Y(n3520));
sg13g2_nand2_2 U4809 (.A(n4323), .B(data_o_6_), .Y(n626));
sg13g2_nor2_2 U4810 (.A(net25928), .B(N1614), .Y(n3684));
sg13g2_nand2_2 U4811 (.A(n3706), .B(n3707), .Y(n4178));
sg13g2_inv_4 U4812 (.A(n4178), .Y(n1775));
sg13g2_nand2_2 U4813 (.A(n4322), .B(data_o_69_), .Y(n628));
sg13g2_o21ai_1 U4814 (.A1(net44327), .A2(three_1), .B1(n4265), .Y(r372_n17));
sg13g2_nand2_2 U4816 (.A(n4323), .B(data_o_88_), .Y(n586));
sg13g2_nor2_2 U4817 (.A(n1134), .B(n168), .Y(n1913));
sg13g2_nor2_2 U4818 (.A(n4333), .B(n3520), .Y(n2244));
sg13g2_nor2_2 U4819 (.A(two_1), .B(N1600), .Y(n3676));
sg13g2_nand2_2 U4820 (.A(n4322), .B(data_o_77_), .Y(n610));
sg13g2_nand2_2 U4821 (.A(n4323), .B(data_o_8_), .Y(n582));
sg13g2_nor2_2 U4822 (.A(addroundkey_round_1), .B(addroundkey_round_2), .Y(net44472));
sg13g2_nand2_2 U4823 (.A(n1905), .B(N1559), .Y(keysched_start_i));
sg13g2_o21ai_1 U4824 (.A1(N1602), .A2(decrypt_i), .B1(n3715), .Y(N313));
sg13g2_o21ai_1 U4825 (.A1(n4242), .A2(n4150), .B1(n4240), .Y(three_3));
sg13g2_nand2_2 U4826 (.A(n4322), .B(data_o_72_), .Y(n620));
sg13g2_nand2_2 U4827 (.A(n4323), .B(data_o_48_), .Y(n674));
sg13g2_inv_4 U4828 (.A(N587), .Y(n3525));
sg13g2_nand2_2 U4829 (.A(net39218), .B(net24695), .Y(net44483));
sg13g2_o21ai_1 U4830 (.A1(N29), .A2(state), .B1(n839), .Y(next_round_2));
sg13g2_nand2_2 U4831 (.A(net47628), .B(n4148), .Y(n4151));
sg13g2_nand2_2 U4832 (.A(n4323), .B(data_o_82_), .Y(n598));
sg13g2_nand2_2 U4833 (.A(n4322), .B(data_o_122_), .Y(n764));
sg13g2_nand3_1 U4834 (.A(addroundkey_ready_o), .B(decrypt_i), .C(N1593), .Y(n3706));
sg13g2_a21oi_2 U4835 (.A1(n2253), .A2(data_i_37_), .B1(n2944), .Y(n2943));
sg13g2_xnor2_1 U4836 (.A(key_i_172_), .B(addroundkey_data_i_108), .Y(n4179));
sg13g2_inv_4 U4837 (.A(n4179), .Y(N749));
sg13g2_nor2_2 U4838 (.A(net44332), .B(n1122), .Y(n1124));
sg13g2_xnor2_1 U4839 (.A(addroundkey_round_0), .B(addroundkey_round_1), .Y(n4273));
sg13g2_o21ai_1 U4840 (.A1(N29), .A2(state), .B1(n834), .Y(next_round_3));
sg13g2_mux2_2 U4841 (.A0(next_last_key_half_62), .A1(last_key_half_62), .S(net24419), .X(n4029));
sg13g2_nand2_2 U4843 (.A(n4322), .B(data_o_68_), .Y(n630));
sg13g2_inv_4 U4844 (.A(n4324), .Y(n4322));
sg13g2_nand2_2 U4845 (.A(n4323), .B(data_o_9_), .Y(n559));
sg13g2_nand3_1 U4846 (.A(net44340), .B(net26619), .C(n4255), .Y(n4254));
sg13g2_nand2_2 U4847 (.A(N1623), .B(N1627), .Y(n3702));
sg13g2_inv_4 U4848 (.A(n3689), .Y(N1623));
sg13g2_inv_4 U4849 (.A(n3693), .Y(N1627));
sg13g2_o21ai_1 U4850 (.A1(n3705), .A2(N1593), .B1(n3708), .Y(n4181));
sg13g2_inv_4 U4851 (.A(n4181), .Y(n557));
sg13g2_xnor2_1 U4852 (.A(key_i_179_), .B(addroundkey_data_i_115), .Y(n4182));
sg13g2_inv_4 U4853 (.A(n4182), .Y(N742));
sg13g2_o21ai_1 U4854 (.A1(n3175), .A2(state), .B1(n3176), .Y(addroundkey_data_i_15));
sg13g2_o21ai_1 U4855 (.A1(n3105), .A2(state), .B1(n3106), .Y(addroundkey_data_i_21));
sg13g2_o21ai_1 U4856 (.A1(n3095), .A2(state), .B1(n3096), .Y(addroundkey_data_i_22));
sg13g2_o21ai_1 U4857 (.A1(n3085), .A2(state), .B1(n3086), .Y(addroundkey_data_i_23));
sg13g2_o21ai_1 U4858 (.A1(n3075), .A2(state), .B1(n3076), .Y(addroundkey_data_i_24));
sg13g2_o21ai_1 U4859 (.A1(n3025), .A2(state), .B1(n3026), .Y(addroundkey_data_i_29));
sg13g2_o21ai_1 U4860 (.A1(n2935), .A2(state), .B1(n2936), .Y(addroundkey_data_i_37));
sg13g2_o21ai_1 U4861 (.A1(n2795), .A2(state), .B1(n2796), .Y(addroundkey_data_i_4));
sg13g2_o21ai_1 U4862 (.A1(n2465), .A2(state), .B1(n2466), .Y(addroundkey_data_i_7));
sg13g2_nor2_2 U4863 (.A(net44327), .B(n1122), .Y(n1126));
sg13g2_mux2_2 U4864 (.A0(next_last_key_half_28), .A1(last_key_half_28), .S(net24419), .X(n3972));
sg13g2_nand2_2 U4866 (.A(r371_n27), .B(n847), .Y(n845));
sg13g2_nand2_2 U4867 (.A(net47628), .B(net47612), .Y(net47660));
sg13g2_xnor2_1 U4868 (.A(net25972), .B(addroundkey_round_0), .Y(r373_n19));
sg13g2_o21ai_1 U4869 (.A1(net44340), .A2(three_3), .B1(n4292), .Y(n4294));
sg13g2_a21oi_2 U4870 (.A1(N29), .A2(addroundkey_ready_o), .B1(n4184), .Y(n3708));
sg13g2_inv_4 U4871 (.A(n3710), .Y(n4184));
sg13g2_o21ai_1 U4872 (.A1(net24787), .A2(n1010), .B1(n2027), .Y(keysched_last_key_i_31));
sg13g2_xnor2_1 U4873 (.A(key_i_168_), .B(addroundkey_data_i_104), .Y(n4185));
sg13g2_inv_4 U4874 (.A(n4185), .Y(N753));
sg13g2_xnor2_1 U4875 (.A(key_i_169_), .B(addroundkey_data_i_105), .Y(n4186));
sg13g2_inv_4 U4876 (.A(n4186), .Y(N752));
sg13g2_xnor2_1 U4877 (.A(key_i_170_), .B(addroundkey_data_i_106), .Y(n4187));
sg13g2_inv_4 U4878 (.A(n4187), .Y(N751));
sg13g2_xnor2_1 U4879 (.A(key_i_171_), .B(addroundkey_data_i_107), .Y(n4188));
sg13g2_inv_4 U4880 (.A(n4188), .Y(N750));
sg13g2_xnor2_1 U4881 (.A(key_i_173_), .B(addroundkey_data_i_109), .Y(n4189));
sg13g2_inv_4 U4882 (.A(n4189), .Y(N748));
sg13g2_xnor2_1 U4883 (.A(key_i_74_), .B(addroundkey_data_i_10), .Y(n4190));
sg13g2_inv_4 U4884 (.A(n4190), .Y(N847));
sg13g2_xnor2_1 U4885 (.A(key_i_174_), .B(addroundkey_data_i_110), .Y(n4191));
sg13g2_inv_4 U4886 (.A(n4191), .Y(N747));
sg13g2_xnor2_1 U4887 (.A(key_i_175_), .B(addroundkey_data_i_111), .Y(n4192));
sg13g2_inv_4 U4888 (.A(n4192), .Y(N746));
sg13g2_xnor2_1 U4889 (.A(key_i_176_), .B(addroundkey_data_i_112), .Y(n4193));
sg13g2_inv_4 U4890 (.A(n4193), .Y(N745));
sg13g2_xnor2_1 U4891 (.A(key_i_177_), .B(addroundkey_data_i_113), .Y(n4194));
sg13g2_inv_4 U4892 (.A(n4194), .Y(N744));
sg13g2_xnor2_1 U4893 (.A(key_i_178_), .B(addroundkey_data_i_114), .Y(n4195));
sg13g2_inv_4 U4894 (.A(n4195), .Y(N743));
sg13g2_xnor2_1 U4895 (.A(key_i_180_), .B(addroundkey_data_i_116), .Y(n4196));
sg13g2_inv_4 U4896 (.A(n4196), .Y(N741));
sg13g2_xnor2_1 U4897 (.A(key_i_181_), .B(addroundkey_data_i_117), .Y(n4197));
sg13g2_inv_4 U4898 (.A(n4197), .Y(N740));
sg13g2_xnor2_1 U4899 (.A(key_i_182_), .B(addroundkey_data_i_118), .Y(n4198));
sg13g2_inv_4 U4900 (.A(n4198), .Y(N739));
sg13g2_xnor2_1 U4901 (.A(key_i_183_), .B(addroundkey_data_i_119), .Y(n4199));
sg13g2_inv_4 U4902 (.A(n4199), .Y(N738));
sg13g2_xnor2_1 U4903 (.A(key_i_75_), .B(addroundkey_data_i_11), .Y(n4200));
sg13g2_inv_4 U4904 (.A(n4200), .Y(N846));
sg13g2_xnor2_1 U4905 (.A(key_i_184_), .B(addroundkey_data_i_120), .Y(n4201));
sg13g2_inv_4 U4906 (.A(n4201), .Y(N737));
sg13g2_xnor2_1 U4907 (.A(key_i_185_), .B(addroundkey_data_i_121), .Y(n4202));
sg13g2_inv_4 U4908 (.A(n4202), .Y(N736));
sg13g2_xnor2_1 U4909 (.A(key_i_186_), .B(addroundkey_data_i_122), .Y(n4203));
sg13g2_inv_4 U4910 (.A(n4203), .Y(N735));
sg13g2_xnor2_1 U4911 (.A(key_i_187_), .B(addroundkey_data_i_123), .Y(n4204));
sg13g2_inv_4 U4912 (.A(n4204), .Y(N734));
sg13g2_o21ai_1 U4913 (.A1(n3245), .A2(state), .B1(n3246), .Y(addroundkey_data_i_124));
sg13g2_o21ai_1 U4914 (.A1(n3235), .A2(state), .B1(n3236), .Y(addroundkey_data_i_125));
sg13g2_o21ai_1 U4915 (.A1(n3225), .A2(state), .B1(n3226), .Y(addroundkey_data_i_126));
sg13g2_o21ai_1 U4916 (.A1(n3215), .A2(state), .B1(n3216), .Y(addroundkey_data_i_127));
sg13g2_o21ai_1 U4917 (.A1(n3205), .A2(state), .B1(n3206), .Y(addroundkey_data_i_12));
sg13g2_o21ai_1 U4918 (.A1(n3195), .A2(state), .B1(n3196), .Y(addroundkey_data_i_13));
sg13g2_o21ai_1 U4919 (.A1(n3185), .A2(state), .B1(n3186), .Y(addroundkey_data_i_14));
sg13g2_o21ai_1 U4920 (.A1(n3165), .A2(state), .B1(n3166), .Y(addroundkey_data_i_16));
sg13g2_o21ai_1 U4921 (.A1(n3155), .A2(state), .B1(n3156), .Y(addroundkey_data_i_17));
sg13g2_o21ai_1 U4922 (.A1(n3135), .A2(state), .B1(n3136), .Y(addroundkey_data_i_19));
sg13g2_o21ai_1 U4923 (.A1(n3125), .A2(state), .B1(n3126), .Y(addroundkey_data_i_1));
sg13g2_o21ai_1 U4924 (.A1(n3115), .A2(state), .B1(n3116), .Y(addroundkey_data_i_20));
sg13g2_o21ai_1 U4925 (.A1(n3065), .A2(state), .B1(n3066), .Y(addroundkey_data_i_25));
sg13g2_o21ai_1 U4926 (.A1(n3055), .A2(state), .B1(n3056), .Y(addroundkey_data_i_26));
sg13g2_o21ai_1 U4927 (.A1(n3045), .A2(state), .B1(n3046), .Y(addroundkey_data_i_27));
sg13g2_o21ai_1 U4928 (.A1(n3035), .A2(state), .B1(n3036), .Y(addroundkey_data_i_28));
sg13g2_o21ai_1 U4929 (.A1(n3015), .A2(state), .B1(n3016), .Y(addroundkey_data_i_2));
sg13g2_o21ai_1 U4930 (.A1(n3005), .A2(state), .B1(n3006), .Y(addroundkey_data_i_30));
sg13g2_o21ai_1 U4931 (.A1(n2995), .A2(state), .B1(n2996), .Y(addroundkey_data_i_31));
sg13g2_o21ai_1 U4932 (.A1(n2985), .A2(state), .B1(n2986), .Y(addroundkey_data_i_32));
sg13g2_o21ai_1 U4933 (.A1(n2975), .A2(state), .B1(n2976), .Y(addroundkey_data_i_33));
sg13g2_o21ai_1 U4934 (.A1(n2965), .A2(state), .B1(n2966), .Y(addroundkey_data_i_34));
sg13g2_o21ai_1 U4935 (.A1(n2955), .A2(state), .B1(n2956), .Y(addroundkey_data_i_35));
sg13g2_o21ai_1 U4936 (.A1(n2945), .A2(state), .B1(n2946), .Y(addroundkey_data_i_36));
sg13g2_o21ai_1 U4937 (.A1(n2925), .A2(state), .B1(n2926), .Y(addroundkey_data_i_38));
sg13g2_o21ai_1 U4938 (.A1(n2915), .A2(state), .B1(n2916), .Y(addroundkey_data_i_39));
sg13g2_o21ai_1 U4939 (.A1(n2905), .A2(state), .B1(n2906), .Y(addroundkey_data_i_3));
sg13g2_o21ai_1 U4940 (.A1(n2895), .A2(state), .B1(n2896), .Y(addroundkey_data_i_40));
sg13g2_o21ai_1 U4941 (.A1(n2885), .A2(state), .B1(n2886), .Y(addroundkey_data_i_41));
sg13g2_o21ai_1 U4942 (.A1(n2875), .A2(state), .B1(n2876), .Y(addroundkey_data_i_42));
sg13g2_o21ai_1 U4943 (.A1(n2865), .A2(state), .B1(n2866), .Y(addroundkey_data_i_43));
sg13g2_o21ai_1 U4944 (.A1(n2855), .A2(state), .B1(n2856), .Y(addroundkey_data_i_44));
sg13g2_o21ai_1 U4945 (.A1(n2845), .A2(state), .B1(n2846), .Y(addroundkey_data_i_45));
sg13g2_o21ai_1 U4946 (.A1(n2835), .A2(state), .B1(n2836), .Y(addroundkey_data_i_46));
sg13g2_o21ai_1 U4947 (.A1(n2815), .A2(state), .B1(n2816), .Y(addroundkey_data_i_48));
sg13g2_o21ai_1 U4948 (.A1(n2805), .A2(state), .B1(n2806), .Y(addroundkey_data_i_49));
sg13g2_o21ai_1 U4949 (.A1(n2785), .A2(state), .B1(n2786), .Y(addroundkey_data_i_50));
sg13g2_o21ai_1 U4950 (.A1(n2775), .A2(state), .B1(n2776), .Y(addroundkey_data_i_51));
sg13g2_o21ai_1 U4951 (.A1(n2765), .A2(state), .B1(n2766), .Y(addroundkey_data_i_52));
sg13g2_o21ai_1 U4952 (.A1(n2755), .A2(state), .B1(n2756), .Y(addroundkey_data_i_53));
sg13g2_o21ai_1 U4953 (.A1(n2745), .A2(state), .B1(n2746), .Y(addroundkey_data_i_54));
sg13g2_o21ai_1 U4954 (.A1(n2735), .A2(state), .B1(n2736), .Y(addroundkey_data_i_55));
sg13g2_o21ai_1 U4955 (.A1(n2725), .A2(state), .B1(n2726), .Y(addroundkey_data_i_56));
sg13g2_o21ai_1 U4956 (.A1(n2715), .A2(state), .B1(n2716), .Y(addroundkey_data_i_57));
sg13g2_o21ai_1 U4957 (.A1(n2705), .A2(state), .B1(n2706), .Y(addroundkey_data_i_58));
sg13g2_o21ai_1 U4958 (.A1(n2695), .A2(state), .B1(n2696), .Y(addroundkey_data_i_59));
sg13g2_o21ai_1 U4959 (.A1(n2685), .A2(state), .B1(n2686), .Y(addroundkey_data_i_5));
sg13g2_o21ai_1 U4960 (.A1(n2675), .A2(state), .B1(n2676), .Y(addroundkey_data_i_60));
sg13g2_o21ai_1 U4961 (.A1(n2665), .A2(state), .B1(n2666), .Y(addroundkey_data_i_61));
sg13g2_o21ai_1 U4962 (.A1(n2655), .A2(state), .B1(n2656), .Y(addroundkey_data_i_62));
sg13g2_o21ai_1 U4963 (.A1(n2645), .A2(state), .B1(n2646), .Y(addroundkey_data_i_63));
sg13g2_o21ai_1 U4964 (.A1(n2635), .A2(state), .B1(n2636), .Y(addroundkey_data_i_64));
sg13g2_o21ai_1 U4965 (.A1(n2625), .A2(state), .B1(n2626), .Y(addroundkey_data_i_65));
sg13g2_o21ai_1 U4966 (.A1(n2615), .A2(state), .B1(n2616), .Y(addroundkey_data_i_66));
sg13g2_o21ai_1 U4967 (.A1(n2605), .A2(state), .B1(n2606), .Y(addroundkey_data_i_67));
sg13g2_o21ai_1 U4968 (.A1(n2595), .A2(state), .B1(n2596), .Y(addroundkey_data_i_68));
sg13g2_o21ai_1 U4969 (.A1(n2575), .A2(state), .B1(n2576), .Y(addroundkey_data_i_6));
sg13g2_o21ai_1 U4970 (.A1(n2565), .A2(state), .B1(n2566), .Y(addroundkey_data_i_70));
sg13g2_o21ai_1 U4971 (.A1(n2555), .A2(state), .B1(n2556), .Y(addroundkey_data_i_71));
sg13g2_o21ai_1 U4972 (.A1(n2545), .A2(state), .B1(n2546), .Y(addroundkey_data_i_72));
sg13g2_o21ai_1 U4973 (.A1(n2525), .A2(state), .B1(n2526), .Y(addroundkey_data_i_74));
sg13g2_o21ai_1 U4974 (.A1(n2515), .A2(state), .B1(n2516), .Y(addroundkey_data_i_75));
sg13g2_o21ai_1 U4975 (.A1(n2505), .A2(state), .B1(n2506), .Y(addroundkey_data_i_76));
sg13g2_o21ai_1 U4976 (.A1(n2495), .A2(state), .B1(n2496), .Y(addroundkey_data_i_77));
sg13g2_o21ai_1 U4977 (.A1(n2485), .A2(state), .B1(n2486), .Y(addroundkey_data_i_78));
sg13g2_o21ai_1 U4978 (.A1(n2475), .A2(state), .B1(n2476), .Y(addroundkey_data_i_79));
sg13g2_o21ai_1 U4979 (.A1(n2455), .A2(state), .B1(n2456), .Y(addroundkey_data_i_80));
sg13g2_o21ai_1 U4980 (.A1(n2445), .A2(state), .B1(n2446), .Y(addroundkey_data_i_81));
sg13g2_o21ai_1 U4981 (.A1(n2435), .A2(state), .B1(n2436), .Y(addroundkey_data_i_82));
sg13g2_o21ai_1 U4982 (.A1(n2425), .A2(state), .B1(n2426), .Y(addroundkey_data_i_83));
sg13g2_o21ai_1 U4983 (.A1(n2415), .A2(state), .B1(n2416), .Y(addroundkey_data_i_84));
sg13g2_o21ai_1 U4984 (.A1(n2405), .A2(state), .B1(n2406), .Y(addroundkey_data_i_85));
sg13g2_o21ai_1 U4985 (.A1(n2395), .A2(state), .B1(n2396), .Y(addroundkey_data_i_86));
sg13g2_o21ai_1 U4986 (.A1(n2385), .A2(state), .B1(n2386), .Y(addroundkey_data_i_87));
sg13g2_o21ai_1 U4987 (.A1(n2375), .A2(state), .B1(n2376), .Y(addroundkey_data_i_88));
sg13g2_o21ai_1 U4988 (.A1(n2365), .A2(state), .B1(n2366), .Y(addroundkey_data_i_89));
sg13g2_o21ai_1 U4989 (.A1(n2355), .A2(state), .B1(n2356), .Y(addroundkey_data_i_8));
sg13g2_o21ai_1 U4990 (.A1(n2345), .A2(state), .B1(n2346), .Y(addroundkey_data_i_90));
sg13g2_o21ai_1 U4991 (.A1(n2335), .A2(state), .B1(n2336), .Y(addroundkey_data_i_91));
sg13g2_o21ai_1 U4992 (.A1(n2325), .A2(state), .B1(n2326), .Y(addroundkey_data_i_92));
sg13g2_o21ai_1 U4993 (.A1(n2315), .A2(state), .B1(n2316), .Y(addroundkey_data_i_93));
sg13g2_o21ai_1 U4994 (.A1(n2305), .A2(state), .B1(n2306), .Y(addroundkey_data_i_94));
sg13g2_o21ai_1 U4995 (.A1(n2295), .A2(state), .B1(n2296), .Y(addroundkey_data_i_95));
sg13g2_o21ai_1 U4996 (.A1(n2285), .A2(state), .B1(n2286), .Y(addroundkey_data_i_96));
sg13g2_o21ai_1 U4997 (.A1(n2275), .A2(state), .B1(n2276), .Y(addroundkey_data_i_97));
sg13g2_o21ai_1 U4998 (.A1(n2265), .A2(state), .B1(n2266), .Y(addroundkey_data_i_98));
sg13g2_o21ai_1 U4999 (.A1(n2255), .A2(state), .B1(n2256), .Y(addroundkey_data_i_99));
sg13g2_o21ai_1 U5000 (.A1(n2242), .A2(state), .B1(n2243), .Y(addroundkey_data_i_9));
sg13g2_a21oi_2 U5001 (.A1(n1120), .A2(N1536), .B1(n1126), .Y(n4205));
sg13g2_inv_4 U5002 (.A(n4205), .Y(next_addroundkey_round_1));
sg13g2_inv_4 U5003 (.A(n4273), .Y(N1536));
sg13g2_mux2_2 U5004 (.A0(next_addroundkey_data_reg_73), .A1(data_o_73_), .S(net24419), .X(n4055));
sg13g2_o21ai_1 U5006 (.A1(n1115), .A2(state), .B1(n1116), .Y(next_addroundkey_start_i));
sg13g2_nor2_2 U5007 (.A(n4217), .B(net26020), .Y(n4207));
sg13g2_inv_4 U5008 (.A(net44483), .Y(net44474));
sg13g2_inv_4 U5009 (.A(net47651), .Y(net47654));
sg13g2_inv_4 U5010 (.A(N1614), .Y(n3683));
sg13g2_nand2_2 U5011 (.A(net47628), .B(N1), .Y(N1614));
sg13g2_nand2_2 U5012 (.A(n3728), .B(n3734), .Y(net39403));
sg13g2_nor2_2 U5013 (.A(r373_n17), .B(r373_n15), .Y(r373_n13));
sg13g2_nand2_2 U5014 (.A(net27521), .B(two_2), .Y(n4146));
sg13g2_nand2_2 U5015 (.A(N1645), .B(keysched_ready_o), .Y(net27301));
sg13g2_inv_4 U5016 (.A(N1657), .Y(n3728));
sg13g2_xnor2_1 U5017 (.A(net47703), .B(n4149), .Y(three_2));
sg13g2_nand2_2 U5018 (.A(keysched_new_key_o_10), .B(net24851), .Y(n2214));
sg13g2_nor2_2 U5019 (.A(r371_n10), .B(r371_n12), .Y(n4208));
sg13g2_nand2_2 U5020 (.A(n3722), .B(n3727), .Y(n4209));
sg13g2_inv_4 U5021 (.A(two_1), .Y(r371_n27));
sg13g2_nand2_2 U5022 (.A(keysched_new_key_o_19), .B(n4156), .Y(n2041));
sg13g2_inv_4 U5023 (.A(n4220), .Y(n4221));
sg13g2_inv_4 U5024 (.A(net24823), .Y(net26188));
sg13g2_inv_4 U5025 (.A(net24783), .Y(n4220));
sg13g2_nand2_2 U5026 (.A(three_0), .B(n3684), .Y(N1620));
sg13g2_inv_4 U5027 (.A(net24419), .Y(net24415));
sg13g2_inv_4 U5028 (.A(n2253), .Y(n4309));
sg13g2_inv_4 U5029 (.A(n4309), .Y(n4307));
sg13g2_nand2_2 U5030 (.A(N7), .B(n3681), .Y(N1571));
sg13g2_inv_4 U5031 (.A(n4214), .Y(n4230));
sg13g2_inv_4 U5032 (.A(net26049), .Y(net25895));
sg13g2_nand2_2 U5033 (.A(net39403), .B(keysched_ready_o), .Y(n4210));
sg13g2_inv_4 U5034 (.A(n3702), .Y(N1118));
sg13g2_o21ai_1 U5035 (.A1(n866), .A2(net24827), .B1(n1979), .Y(keysched_last_key_i_6));
sg13g2_nand2_2 U5036 (.A(net26529), .B(subbytes_sbox_data_o_6), .Y(net26531));
sg13g2_o21ai_1 U5037 (.A1(net24795), .A2(n2095), .B1(n2096), .Y(keysched_last_key_i_166));
sg13g2_o21ai_1 U5038 (.A1(net26188), .A2(n2147), .B1(n2148), .Y(keysched_last_key_i_141));
sg13g2_o21ai_1 U5039 (.A1(n4211), .A2(n1054), .B1(n2038), .Y(keysched_last_key_i_21));
sg13g2_o21ai_1 U5040 (.A1(net24791), .A2(n2072), .B1(n2073), .Y(keysched_last_key_i_177));
sg13g2_o21ai_1 U5041 (.A1(net24791), .A2(n2068), .B1(n2069), .Y(keysched_last_key_i_179));
sg13g2_inv_4 U5042 (.A(n4175), .Y(net39311));
sg13g2_o21ai_1 U5043 (.A1(n4221), .A2(n2139), .B1(n2140), .Y(keysched_last_key_i_145));
sg13g2_o21ai_1 U5044 (.A1(net26210), .A2(n930), .B1(n2007), .Y(keysched_last_key_i_4));
sg13g2_o21ai_1 U5045 (.A1(net24801), .A2(n1046), .B1(n2036), .Y(keysched_last_key_i_23));
sg13g2_inv_4 U5046 (.A(net44320), .Y(next_addroundkey_ready_o));
sg13g2_nand2_2 U5047 (.A(net44482), .B(net44483), .Y(net44320));
sg13g2_nand2_2 U5048 (.A(n3733), .B(n3729), .Y(N1657));
sg13g2_inv_4 U5049 (.A(net24821), .Y(net24783));
sg13g2_inv_4 U5050 (.A(n1905), .Y(n4212));
sg13g2_o21ai_1 U5051 (.A1(net24795), .A2(n2042), .B1(n2043), .Y(keysched_last_key_i_191));
sg13g2_o21ai_1 U5052 (.A1(net24795), .A2(n2093), .B1(n2094), .Y(keysched_last_key_i_167));
sg13g2_o21ai_1 U5053 (.A1(net24787), .A2(n1050), .B1(n2037), .Y(keysched_last_key_i_22));
sg13g2_inv_4 U5054 (.A(net24821), .Y(net24787));
sg13g2_nand2_2 U5055 (.A(N1645), .B(keysched_ready_o), .Y(n4214));
sg13g2_inv_4 U5056 (.A(net24875), .Y(net24837));
sg13g2_nand2_2 U5057 (.A(three_3), .B(net44340), .Y(n4292));
sg13g2_nor2_2 U5058 (.A(net47703), .B(n4149), .Y(n4150));
sg13g2_inv_4 U5059 (.A(net25885), .Y(net24847));
sg13g2_nand2_2 U5060 (.A(net26947), .B(n4219), .Y(n4217));
sg13g2_nor2_2 U5061 (.A(net39212), .B(n4277), .Y(n4279));
sg13g2_o21ai_1 U5062 (.A1(n4332), .A2(n3395), .B1(n3396), .Y(addroundkey_data_i_110));
sg13g2_o21ai_1 U5063 (.A1(n4332), .A2(n3325), .B1(n3326), .Y(addroundkey_data_i_117));
sg13g2_o21ai_1 U5064 (.A1(n4332), .A2(n3335), .B1(n3336), .Y(addroundkey_data_i_116));
sg13g2_o21ai_1 U5065 (.A1(n4332), .A2(n3355), .B1(n3356), .Y(addroundkey_data_i_114));
sg13g2_o21ai_1 U5066 (.A1(n4332), .A2(n3375), .B1(n3376), .Y(addroundkey_data_i_112));
sg13g2_o21ai_1 U5067 (.A1(n4332), .A2(n3445), .B1(n3446), .Y(addroundkey_data_i_106));
sg13g2_inv_4 U5068 (.A(n4331), .Y(n4332));
sg13g2_nand2_2 U5069 (.A(subbytes_ready_o), .B(N313), .Y(n843));
sg13g2_nand2_2 U5070 (.A(n3716), .B(n3721), .Y(n4218));
sg13g2_o21ai_1 U5071 (.A1(net24791), .A2(n2082), .B1(n2083), .Y(keysched_last_key_i_172));
sg13g2_o21ai_1 U5072 (.A1(net24791), .A2(n2076), .B1(n2077), .Y(keysched_last_key_i_175));
sg13g2_o21ai_1 U5073 (.A1(net24791), .A2(n2047), .B1(n2048), .Y(keysched_last_key_i_189));
sg13g2_nand2_2 U5074 (.A(net24881), .B(keysched_new_key_o_6), .Y(n1979));
sg13g2_inv_4 U5075 (.A(net27680), .Y(net24863));
sg13g2_nand2_2 U5076 (.A(keysched_new_key_o_14), .B(n4239), .Y(n2130));
sg13g2_inv_4 U5077 (.A(n560), .Y(n4324));
sg13g2_inv_4 U5078 (.A(n4324), .Y(n4320));
sg13g2_inv_4 U5079 (.A(n4314), .Y(n4312));
sg13g2_nand2_2 U5080 (.A(net38935), .B(n4230), .Y(n4281));
sg13g2_inv_4 U5081 (.A(n4162), .Y(n4293));
sg13g2_inv_4 U5082 (.A(n4311), .Y(n4310));
sg13g2_inv_4 U5083 (.A(n4295), .Y(n4298));
sg13g2_nand2_2 U5084 (.A(net39311), .B(net43702), .Y(n4278));
sg13g2_inv_4 U5085 (.A(net24633), .Y(net24601));
sg13g2_inv_4 U5086 (.A(net47628), .Y(net26538));
sg13g2_nand2_2 U5087 (.A(net26019), .B(net44816), .Y(net44819));
sg13g2_inv_4 U5088 (.A(state), .Y(n4333));
sg13g2_inv_4 U5090 (.A(n4314), .Y(n4313));
sg13g2_inv_4 U5091 (.A(n4275), .Y(n4276));
sg13g2_inv_4 U5092 (.A(sbox_data_o_0), .Y(n4275));
sg13g2_inv_4 U5093 (.A(sbox_data_o_3), .Y(n4288));
sg13g2_inv_4 U5094 (.A(n4288), .Y(n4289));
sg13g2_inv_4 U5095 (.A(net24875), .Y(net25892));
sg13g2_inv_4 U5096 (.A(n4309), .Y(n4308));
sg13g2_inv_4 U5097 (.A(n2244), .Y(n4314));
sg13g2_inv_4 U5098 (.A(net24419), .Y(net24383));
sg13g2_inv_4 U5099 (.A(net24419), .Y(net24381));
sg13g2_inv_4 U5100 (.A(net24419), .Y(net24393));
sg13g2_inv_4 U5103 (.A(net25928), .Y(two_1));
sg13g2_inv_4 U5104 (.A(n1913), .Y(N1559));
sg13g2_inv_4 U5105 (.A(n851), .Y(n4315));
sg13g2_inv_4 U5106 (.A(n1134), .Y(net38935));
sg13g2_inv_4 U5109 (.A(n4283), .Y(net24743));
sg13g2_inv_4 U5110 (.A(N1559), .Y(net24419));
sg13g2_inv_4 U5111 (.A(keysched_sbox_access_o), .Y(n4252));
sg13g2_o21ai_1 U5112 (.A1(n4211), .A2(n1074), .B1(n2067), .Y(keysched_last_key_i_17));
sg13g2_inv_4 U5113 (.A(key_i_15_), .Y(n1082));
sg13g2_nand2_2 U5114 (.A(n4209), .B(keysched_ready_o), .Y(n4228));
sg13g2_a21oi_2 U5115 (.A1(n2244), .A2(n3207), .B1(n3208), .Y(n3206));
sg13g2_o21ai_1 U5116 (.A1(net24791), .A2(n2074), .B1(n2075), .Y(keysched_last_key_i_176));
sg13g2_inv_4 U5117 (.A(sbox_data_o_4), .Y(n4222));
sg13g2_inv_4 U5118 (.A(n4222), .Y(n4223));
sg13g2_o21ai_1 U5119 (.A1(n4221), .A2(n966), .B1(n2016), .Y(keysched_last_key_i_41));
sg13g2_o21ai_1 U5120 (.A1(n4221), .A2(n2051), .B1(n2052), .Y(keysched_last_key_i_187));
sg13g2_o21ai_1 U5121 (.A1(n4332), .A2(n3295), .B1(n3296), .Y(addroundkey_data_i_11));
sg13g2_a21oi_2 U5122 (.A1(n4312), .A2(n3327), .B1(n3328), .Y(n3326));
sg13g2_a21oi_2 U5123 (.A1(n4312), .A2(n3337), .B1(n3338), .Y(n3336));
sg13g2_a21oi_2 U5124 (.A1(n4312), .A2(n3347), .B1(n3348), .Y(n3346));
sg13g2_a21oi_2 U5125 (.A1(n4312), .A2(n3357), .B1(n3358), .Y(n3356));
sg13g2_a21oi_2 U5126 (.A1(n4312), .A2(n3377), .B1(n3378), .Y(n3376));
sg13g2_a21oi_2 U5127 (.A1(n4312), .A2(n3387), .B1(n3388), .Y(n3386));
sg13g2_a21oi_2 U5128 (.A1(n4312), .A2(n3367), .B1(n3368), .Y(n3366));
sg13g2_o21ai_1 U5129 (.A1(net24795), .A2(n2055), .B1(n2056), .Y(keysched_last_key_i_185));
sg13g2_o21ai_1 U5130 (.A1(n4221), .A2(n2053), .B1(n2054), .Y(keysched_last_key_i_186));
sg13g2_a21oi_2 U5131 (.A1(n2244), .A2(n3297), .B1(n3298), .Y(n3296));
sg13g2_inv_4 U5132 (.A(n4275), .Y(n4224));
sg13g2_inv_4 U5133 (.A(n4288), .Y(n4225));
sg13g2_o21ai_1 U5134 (.A1(n4332), .A2(n3255), .B1(n3256), .Y(addroundkey_data_i_123));
sg13g2_a21oi_2 U5135 (.A1(n2244), .A2(n3257), .B1(n3258), .Y(n3256));
sg13g2_o21ai_1 U5136 (.A1(n4332), .A2(n3275), .B1(n3276), .Y(addroundkey_data_i_121));
sg13g2_a21oi_2 U5137 (.A1(n4313), .A2(n3277), .B1(n3278), .Y(n3276));
sg13g2_mux2_2 U5138 (.A0(data_o_11_), .A1(next_addroundkey_data_reg_11), .S(net24393), .X(n4117));
sg13g2_o21ai_1 U5139 (.A1(n4332), .A2(n3285), .B1(n3286), .Y(addroundkey_data_i_120));
sg13g2_a21oi_2 U5140 (.A1(n2244), .A2(n3287), .B1(n3288), .Y(n3286));
sg13g2_o21ai_1 U5141 (.A1(n4332), .A2(n3265), .B1(n3266), .Y(addroundkey_data_i_122));
sg13g2_a21oi_2 U5142 (.A1(n4313), .A2(n3267), .B1(n3268), .Y(n3266));
sg13g2_o21ai_1 U5143 (.A1(n4332), .A2(n3305), .B1(n3306), .Y(addroundkey_data_i_119));
sg13g2_a21oi_2 U5144 (.A1(n4313), .A2(n3307), .B1(n3308), .Y(n3306));
sg13g2_o21ai_1 U5145 (.A1(n4332), .A2(n3315), .B1(n3316), .Y(addroundkey_data_i_118));
sg13g2_a21oi_2 U5146 (.A1(n2244), .A2(n3317), .B1(n3318), .Y(n3316));
sg13g2_o21ai_1 U5147 (.A1(net26188), .A2(n1950), .B1(n1951), .Y(keysched_last_key_i_83));
sg13g2_o21ai_1 U5148 (.A1(net26188), .A2(n1952), .B1(n1953), .Y(keysched_last_key_i_82));
sg13g2_o21ai_1 U5149 (.A1(net26188), .A2(n2225), .B1(n2226), .Y(keysched_last_key_i_104));
sg13g2_o21ai_1 U5150 (.A1(net26188), .A2(n2223), .B1(n2224), .Y(keysched_last_key_i_105));
sg13g2_inv_4 U5151 (.A(n4226), .Y(n4227));
sg13g2_a21oi_2 U5152 (.A1(last_key_half_46), .A2(net26864), .B1(n948), .Y(n947));
sg13g2_inv_4 U5153 (.A(net24881), .Y(net27680));
sg13g2_inv_4 U5154 (.A(net25885), .Y(net24849));
sg13g2_inv_4 U5155 (.A(r371_n17), .Y(n4246));
sg13g2_nand2_2 U5156 (.A(net47703), .B(net47653), .Y(N1611));
sg13g2_nand2_2 U5157 (.A(N1324), .B(N1123), .Y(n3734));
sg13g2_o21ai_1 U5158 (.A1(n4221), .A2(n2091), .B1(n2092), .Y(keysched_last_key_i_168));
sg13g2_nand2_2 U5159 (.A(net44483), .B(net44493), .Y(net44768));
sg13g2_inv_4 U5160 (.A(r370_n12), .Y(n4245));
sg13g2_nand2_2 U5161 (.A(state), .B(n3520), .Y(n2248));
sg13g2_o21ai_1 U5162 (.A1(n4332), .A2(n3405), .B1(n3406), .Y(addroundkey_data_i_10));
sg13g2_a21oi_2 U5163 (.A1(n4312), .A2(n3407), .B1(n3408), .Y(n3406));
sg13g2_inv_4 U5164 (.A(n4146), .Y(n4145));
sg13g2_o21ai_1 U5165 (.A1(n4327), .A2(n755), .B1(n756), .Y(subbytes_data_i_126));
sg13g2_nand2_2 U5166 (.A(N29), .B(N1610), .Y(n4229));
sg13g2_inv_4 U5167 (.A(two_2), .Y(r371_n28));
sg13g2_o21ai_1 U5168 (.A1(n4327), .A2(n635), .B1(n636), .Y(subbytes_data_i_65));
sg13g2_nand2_2 U5169 (.A(n4143), .B(net47653), .Y(net26619));
sg13g2_o21ai_1 U5170 (.A1(n4325), .A2(n617), .B1(n618), .Y(subbytes_data_i_73));
sg13g2_nand2_2 U5171 (.A(n4245), .B(n4231), .Y(n4232));
sg13g2_inv_4 U5172 (.A(n3692), .Y(N1626));
sg13g2_nand2_2 U5173 (.A(n3683), .B(N1626), .Y(n3704));
sg13g2_nand2_2 U5174 (.A(N1623), .B(N1626), .Y(n3701));
sg13g2_nand2_2 U5175 (.A(N1622), .B(N1626), .Y(n3697));
sg13g2_nand2_2 U5176 (.A(subbytes_data_o_29), .B(n4321), .Y(n1854));
sg13g2_nand2_2 U5177 (.A(n4208), .B(N1119), .Y(n3719));
sg13g2_nor2_2 U5178 (.A(r370_n10), .B(n3704), .Y(n4231));
sg13g2_nand2_2 U5179 (.A(subbytes_data_o_40), .B(n4319), .Y(n1841));
sg13g2_nand2_2 U5180 (.A(net26529), .B(subbytes_sbox_data_o_7), .Y(n4290));
sg13g2_nand2_2 U5181 (.A(net26529), .B(subbytes_sbox_data_o_5), .Y(n4234));
sg13g2_o21ai_1 U5182 (.A1(n4221), .A2(n878), .B1(n1994), .Y(keysched_last_key_i_61));
sg13g2_nand2_2 U5183 (.A(subbytes_data_o_46), .B(n4320), .Y(n1835));
sg13g2_nand2_2 U5184 (.A(subbytes_data_o_55), .B(n4321), .Y(n1825));
sg13g2_nand2_2 U5185 (.A(subbytes_data_o_103), .B(n4316), .Y(n1899));
sg13g2_nand2_2 U5186 (.A(data_o_91_), .B(n4322), .Y(n578));
sg13g2_o21ai_1 U5187 (.A1(n4221), .A2(n1963), .B1(n1964), .Y(keysched_last_key_i_77));
sg13g2_inv_4 U5188 (.A(n4268), .Y(n4269));
sg13g2_o21ai_1 U5189 (.A1(net24787), .A2(n1030), .B1(n2032), .Y(keysched_last_key_i_27));
sg13g2_o21ai_1 U5190 (.A1(net24787), .A2(n1094), .B1(n2172), .Y(keysched_last_key_i_12));
sg13g2_o21ai_1 U5191 (.A1(n4325), .A2(n1338), .B1(n1816), .Y(mixcol_data_i_63));
sg13g2_nand2_2 U5192 (.A(n4297), .B(n614), .Y(subbytes_data_i_75));
sg13g2_nand2_2 U5193 (.A(n822), .B(n4234), .Y(sbox_data_i_5));
sg13g2_inv_4 U5194 (.A(sbox_data_o_5), .Y(n4236));
sg13g2_inv_4 U5195 (.A(n4236), .Y(n4237));
sg13g2_o21ai_1 U5196 (.A1(net24795), .A2(n950), .B1(n2012), .Y(keysched_last_key_i_45));
sg13g2_inv_4 U5197 (.A(N1611), .Y(n3681));
sg13g2_o21ai_1 U5198 (.A1(n4221), .A2(n2158), .B1(n2159), .Y(keysched_last_key_i_136));
sg13g2_nand2_2 U5199 (.A(net26529), .B(subbytes_sbox_data_o_2), .Y(n4267));
sg13g2_nand2_2 U5200 (.A(net26529), .B(subbytes_sbox_data_o_1), .Y(n4285));
sg13g2_nand2_2 U5201 (.A(n4218), .B(keysched_ready_o), .Y(n4238));
sg13g2_o21ai_1 U5202 (.A1(net24787), .A2(n1066), .B1(n2041), .Y(keysched_last_key_i_19));
sg13g2_o21ai_1 U5203 (.A1(n4330), .A2(n761), .B1(n762), .Y(subbytes_data_i_123));
sg13g2_o21ai_1 U5204 (.A1(n4325), .A2(n787), .B1(n788), .Y(subbytes_data_i_111));
sg13g2_nand2_2 U5205 (.A(data_o_111_), .B(n4316), .Y(n788));
sg13g2_inv_4 U5206 (.A(n168), .Y(net39218));
sg13g2_inv_4 U5207 (.A(n4151), .Y(n4241));
sg13g2_inv_4 U5208 (.A(net47653), .Y(n4242));
sg13g2_nand2_2 U5209 (.A(n4241), .B(n4242), .Y(n4240));
sg13g2_inv_4 U5210 (.A(net27680), .Y(net24851));
sg13g2_nand2_2 U5211 (.A(keysched_new_key_o_8), .B(net24863), .Y(n1937));
sg13g2_inv_4 U5212 (.A(net24829), .Y(net26210));
sg13g2_nand2_2 U5213 (.A(keysched_new_key_o_31), .B(net24847), .Y(n2027));
sg13g2_o21ai_1 U5214 (.A1(net24783), .A2(n1022), .B1(n2030), .Y(keysched_last_key_i_29));
sg13g2_nand2_2 U5215 (.A(net26430), .B(keysched_new_key_o_27), .Y(n2032));
sg13g2_nand2_2 U5216 (.A(keysched_new_key_o_22), .B(n4239), .Y(n2037));
sg13g2_nand2_2 U5217 (.A(net26529), .B(subbytes_sbox_data_o_0), .Y(n4287));
sg13g2_nand4_1 U5218 (.A(r370_n13), .B(r370_n19), .C(n4253), .D(n4254), .Y(n3730));
sg13g2_o21ai_1 U5219 (.A1(net24791), .A2(n1078), .B1(n2088), .Y(keysched_last_key_i_16));
sg13g2_nand2_2 U5220 (.A(keysched_new_key_o_16), .B(net24845), .Y(n2088));
sg13g2_nand2_2 U5221 (.A(net44478), .B(net24695), .Y(net44482));
sg13g2_inv_4 U5222 (.A(three_0), .Y(r370_n26));
sg13g2_xnor2_1 U5223 (.A(four_3_), .B(addroundkey_round_3), .Y(n4243));
sg13g2_inv_4 U5224 (.A(n4243), .Y(r373_n10));
sg13g2_nand3_1 U5225 (.A(n4245), .B(n4244), .C(N1116), .Y(n3718));
sg13g2_inv_4 U5226 (.A(r370_n10), .Y(n4244));
sg13g2_inv_4 U5227 (.A(n3703), .Y(N1116));
sg13g2_a21oi_2 U5228 (.A1(n4264), .A2(N1121), .B1(N1648), .Y(n3722));
sg13g2_inv_4 U5230 (.A(n3688), .Y(N1622));
sg13g2_a21oi_2 U5231 (.A1(n1912), .A2(addroundkey_round_0), .B1(n1913), .Y(n1911));
sg13g2_nand4_1 U5232 (.A(r371_n19), .B(n4246), .C(n4263), .D(n4262), .Y(r371_n12));
sg13g2_a21oi_2 U5233 (.A1(key_i_129_), .A2(n4220), .B1(n4247), .Y(n4248));
sg13g2_inv_4 U5234 (.A(n2174), .Y(n4247));
sg13g2_inv_4 U5235 (.A(n4248), .Y(keysched_last_key_i_129));
sg13g2_inv_4 U5236 (.A(net39135), .Y(net44478));
sg13g2_nand3_1 U5237 (.A(n4302), .B(n4303), .C(addroundkey_round_3), .Y(n4300));
sg13g2_a21oi_2 U5238 (.A1(n4207), .A2(net44475), .B1(n4256), .Y(n1914));
sg13g2_nand2_2 U5239 (.A(net44482), .B(net44769), .Y(n4258));
sg13g2_nand2_2 U5240 (.A(r373_n26), .B(two_1), .Y(n3694));
sg13g2_inv_4 U5241 (.A(net25927), .Y(net25928));
sg13g2_inv_4 U5243 (.A(net25927), .Y(net27520));
sg13g2_nand2_2 U5244 (.A(net25927), .B(net47625), .Y(net27332));
sg13g2_inv_4 U5245 (.A(three_0), .Y(net25972));
sg13g2_inv_4 U5246 (.A(two_0), .Y(three_0));
sg13g2_nand2_2 U5247 (.A(net26538), .B(N1), .Y(n3689));
sg13g2_inv_4 U5248 (.A(net47654), .Y(N1));
sg13g2_inv_4 U5250 (.A(net47651), .Y(net47653));
sg13g2_inv_4 U5251 (.A(round_2_), .Y(net47628));
sg13g2_nor2_2 U5252 (.A(net39218), .B(n4249), .Y(net44475));
sg13g2_nand2_2 U5253 (.A(n4207), .B(n168), .Y(net44319));
sg13g2_inv_4 U5254 (.A(net26019), .Y(net26020));
sg13g2_nand2_2 U5255 (.A(n4250), .B(net44340), .Y(n4249));
sg13g2_nor2_2 U5256 (.A(net44474), .B(n4249), .Y(net44473));
sg13g2_nand2_2 U5257 (.A(net44472), .B(net44340), .Y(net44493));
sg13g2_nor2_2 U5258 (.A(n1122), .B(net44340), .Y(n1121));
sg13g2_nor2_2 U5259 (.A(addroundkey_round_1), .B(addroundkey_round_2), .Y(n4250));
sg13g2_inv_4 U5260 (.A(net26537), .Y(net47703));
sg13g2_inv_4 U5262 (.A(net26537), .Y(net26539));
sg13g2_nand2_2 U5263 (.A(net39126), .B(n166), .Y(net26946));
sg13g2_inv_4 U5264 (.A(net26946), .Y(net26947));
sg13g2_inv_4 U5265 (.A(n4228), .Y(net39214));
sg13g2_nand3_1 U5266 (.A(n4238), .B(net39126), .C(n166), .Y(net39135));
sg13g2_inv_4 U5267 (.A(n3696), .Y(N1124));
sg13g2_nand2_2 U5268 (.A(net25972), .B(net25928), .Y(n3691));
sg13g2_nand2_2 U5269 (.A(net26537), .B(net47653), .Y(n3688));
sg13g2_nand2_2 U5270 (.A(net27145), .B(n4251), .Y(r370_n17));
sg13g2_nor2_2 U5271 (.A(r370_n15), .B(r370_n17), .Y(r370_n13));
sg13g2_nand2_2 U5272 (.A(r370_n27), .B(addroundkey_round_1), .Y(n4251));
sg13g2_inv_4 U5273 (.A(one_1_), .Y(r370_n27));
sg13g2_nand2_2 U5274 (.A(one_1_), .B(net44327), .Y(net27145));
sg13g2_o21ai_1 U5275 (.A1(net27521), .A2(three_0), .B1(net27332), .Y(one_1_));
sg13g2_inv_4 U5276 (.A(net27520), .Y(net27521));
sg13g2_xnor2_1 U5277 (.A(net26539), .B(net27332), .Y(one_2_));
sg13g2_nor2_2 U5278 (.A(two_0), .B(four_1), .Y(net47612));
sg13g2_nand2_2 U5279 (.A(four_1), .B(two_0), .Y(n4148));
sg13g2_xnor2_1 U5281 (.A(round_2_), .B(four_1), .Y(two_2));
sg13g2_inv_4 U5282 (.A(net39403), .Y(net39212));
sg13g2_nand2_2 U5283 (.A(N1323), .B(N1120), .Y(n3733));
sg13g2_inv_4 U5284 (.A(n3700), .Y(N1120));
sg13g2_nand2_2 U5285 (.A(r370_n13), .B(r370_n19), .Y(r370_n12));
sg13g2_xnor2_1 U5286 (.A(net44332), .B(one_2_), .Y(r370_n15));
sg13g2_nand2_2 U5287 (.A(n3730), .B(n3731), .Y(N1653));
sg13g2_nand2_2 U5288 (.A(net25972), .B(two_1), .Y(n3693));
sg13g2_nand2_2 U5289 (.A(keysched_sbox_data_o_6), .B(net26029), .Y(n820));
sg13g2_nand2_2 U5290 (.A(n820), .B(net26531), .Y(sbox_data_i_6));
sg13g2_inv_4 U5291 (.A(n4252), .Y(net26029));
sg13g2_nor2_2 U5292 (.A(n815), .B(keysched_sbox_access_o), .Y(sbox_decrypt_i));
sg13g2_nand2_2 U5293 (.A(net26947), .B(n4219), .Y(n2241));
sg13g2_inv_4 U5294 (.A(n2241), .Y(net44816));
sg13g2_nor2_2 U5295 (.A(keysched_ready_o), .B(n1134), .Y(net26019));
sg13g2_inv_4 U5296 (.A(net24695), .Y(n1134));
sg13g2_nand2_2 U5297 (.A(n4254), .B(n4253), .Y(r370_n10));
sg13g2_nand2_2 U5298 (.A(n4144), .B(addroundkey_round_3), .Y(n4253));
sg13g2_nand2_2 U5299 (.A(net26619), .B(n4255), .Y(n4144));
sg13g2_nand2_2 U5300 (.A(net47660), .B(net26618), .Y(n4255));
sg13g2_inv_4 U5301 (.A(net47654), .Y(net26618));
sg13g2_inv_4 U5302 (.A(n4257), .Y(net24883));
sg13g2_inv_4 U5303 (.A(net24883), .Y(net24879));
sg13g2_inv_4 U5304 (.A(net24883), .Y(net24881));
sg13g2_nand3_1 U5305 (.A(n4259), .B(n4258), .C(n1905), .Y(n4257));
sg13g2_inv_4 U5306 (.A(net44768), .Y(net44769));
sg13g2_nand2_2 U5307 (.A(net44816), .B(net44818), .Y(n4259));
sg13g2_nand2_2 U5308 (.A(n168), .B(net44493), .Y(net44654));
sg13g2_inv_4 U5309 (.A(net24829), .Y(net24827));
sg13g2_inv_4 U5310 (.A(n1914), .Y(net24829));
sg13g2_inv_4 U5311 (.A(net24829), .Y(net24825));
sg13g2_inv_4 U5312 (.A(net24829), .Y(net26302));
sg13g2_inv_4 U5313 (.A(n1134), .Y(net43702));
sg13g2_inv_4 U5314 (.A(sbox_data_o_1), .Y(n4260));
sg13g2_nand2_2 U5315 (.A(three_0), .B(n3682), .Y(N1613));
sg13g2_nand2_2 U5316 (.A(data_o_63_), .B(n4321), .Y(n640));
sg13g2_inv_4 U5317 (.A(n4260), .Y(n4261));
sg13g2_nand2_2 U5318 (.A(r371_n28), .B(addroundkey_round_2), .Y(n4262));
sg13g2_nand2_2 U5319 (.A(net47686), .B(net44332), .Y(n4263));
sg13g2_inv_4 U5320 (.A(r371_n28), .Y(net47686));
sg13g2_nor2_2 U5321 (.A(n4294), .B(r372_n12), .Y(n4264));
sg13g2_nand2_2 U5322 (.A(three_1), .B(net44327), .Y(n4265));
sg13g2_nand2_2 U5323 (.A(subbytes_data_o_21), .B(n4318), .Y(n1862));
sg13g2_nand2_2 U5324 (.A(subbytes_data_o_47), .B(n4320), .Y(n1834));
sg13g2_nand2_2 U5325 (.A(subbytes_data_o_51), .B(n4320), .Y(n1829));
sg13g2_nand2_2 U5326 (.A(subbytes_data_o_53), .B(n4320), .Y(n1827));
sg13g2_nand2_2 U5327 (.A(subbytes_data_o_49), .B(n4320), .Y(n1832));
sg13g2_inv_4 U5328 (.A(net47660), .Y(n4143));
sg13g2_nand2_2 U5329 (.A(subbytes_data_o_61), .B(n4321), .Y(n1818));
sg13g2_o21ai_1 U5330 (.A1(net24783), .A2(n1102), .B1(n2214), .Y(keysched_last_key_i_10));
sg13g2_o21ai_1 U5331 (.A1(net24791), .A2(n2049), .B1(n2050), .Y(keysched_last_key_i_188));
sg13g2_inv_4 U5332 (.A(net26029), .Y(net26529));
sg13g2_nand2_2 U5333 (.A(three_0), .B(n3682), .Y(N1593));
sg13g2_nand2_2 U5334 (.A(data_o_83_), .B(n4317), .Y(n596));
sg13g2_o21ai_1 U5335 (.A1(n4326), .A2(n657), .B1(n658), .Y(subbytes_data_i_55));
sg13g2_o21ai_1 U5336 (.A1(n4221), .A2(n2107), .B1(n2108), .Y(keysched_last_key_i_160));
sg13g2_nand2_2 U5337 (.A(keysched_new_key_o_28), .B(n4156), .Y(n2031));
sg13g2_nand2_2 U5338 (.A(net24881), .B(keysched_new_key_o_3), .Y(n2018));
sg13g2_o21ai_1 U5339 (.A1(addroundkey_round_0), .A2(n4213), .B1(n1911), .Y(keysched_round_i_0));
sg13g2_o21ai_1 U5340 (.A1(net24783), .A2(n852), .B1(n4235), .Y(keysched_last_key_i_9));
sg13g2_nand2_2 U5341 (.A(keysched_new_key_o_12), .B(net24851), .Y(n2172));
sg13g2_nand2_2 U5342 (.A(N1613), .B(decrypt_i), .Y(n4266));
sg13g2_nand2_2 U5343 (.A(n4267), .B(n828), .Y(sbox_data_i_2));
sg13g2_nand2_2 U5344 (.A(keysched_sbox_data_o_2), .B(net26029), .Y(n828));
sg13g2_o21ai_1 U5345 (.A1(n4211), .A2(n1038), .B1(n2034), .Y(keysched_last_key_i_25));
sg13g2_nand2_2 U5346 (.A(keysched_new_key_o_188), .B(n4156), .Y(n2050));
sg13g2_nand2_2 U5347 (.A(keysched_new_key_o_183), .B(net24847), .Y(n2060));
sg13g2_nand2_2 U5348 (.A(keysched_new_key_o_17), .B(net24847), .Y(n2067));
sg13g2_inv_4 U5349 (.A(N1571), .Y(n3682));
sg13g2_nand2_2 U5350 (.A(net44319), .B(net44320), .Y(n1912));
sg13g2_nand2_2 U5351 (.A(keysched_new_key_o_23), .B(net26430), .Y(n2036));
sg13g2_o21ai_1 U5352 (.A1(n4325), .A2(n727), .B1(n728), .Y(subbytes_data_i_23));
sg13g2_xnor2_1 U5353 (.A(three_0), .B(net25928), .Y(three_1));
sg13g2_nand2_2 U5354 (.A(n4270), .B(n2193), .Y(keysched_last_key_i_11));
sg13g2_nand2_2 U5355 (.A(net24879), .B(keysched_new_key_o_0), .Y(n2235));
sg13g2_nand2_2 U5356 (.A(net24879), .B(keysched_new_key_o_5), .Y(n1996));
sg13g2_nand2_2 U5357 (.A(keysched_sbox_data_o_5), .B(net26029), .Y(n822));
sg13g2_o21ai_1 U5358 (.A1(net27141), .A2(net44327), .B1(n1910), .Y(keysched_round_i_1));
sg13g2_o21ai_1 U5359 (.A1(net27141), .A2(net44332), .B1(n1909), .Y(keysched_round_i_2));
sg13g2_nand2_2 U5360 (.A(n1907), .B(n4271), .Y(keysched_round_i_3));
sg13g2_o21ai_1 U5361 (.A1(net24795), .A2(n2065), .B1(n2066), .Y(keysched_last_key_i_180));
sg13g2_o21ai_1 U5362 (.A1(n886), .A2(net24825), .B1(n1996), .Y(keysched_last_key_i_5));
sg13g2_nand2_2 U5363 (.A(keysched_new_key_o_29), .B(net24851), .Y(n2030));
sg13g2_nand2_2 U5364 (.A(keysched_new_key_o_15), .B(net24849), .Y(n2109));
sg13g2_nand2_2 U5365 (.A(keysched_new_key_o_20), .B(net24857), .Y(n2039));
sg13g2_nand2_2 U5366 (.A(net24881), .B(keysched_new_key_o_7), .Y(n1958));
sg13g2_buf_8 U5367 (.A(sbox_data_o_6), .X(n4274));
sg13g2_o21ai_1 U5368 (.A1(net24791), .A2(n1070), .B1(n2046), .Y(keysched_last_key_i_18));
sg13g2_inv_4 U5369 (.A(net25885), .Y(net24857));
sg13g2_nand2_2 U5370 (.A(keysched_new_key_o_2), .B(n4156), .Y(n2029));
sg13g2_o21ai_1 U5371 (.A1(n4211), .A2(n1014), .B1(n2028), .Y(keysched_last_key_i_30));
sg13g2_nand2_2 U5372 (.A(n4233), .B(key_i_15_), .Y(n4286));
sg13g2_nand3_1 U5373 (.A(net39214), .B(n4214), .C(net38935), .Y(n4283));
sg13g2_inv_4 U5374 (.A(net24879), .Y(net25885));
sg13g2_o21ai_1 U5375 (.A1(net24787), .A2(n1086), .B1(n2130), .Y(keysched_last_key_i_14));
sg13g2_nand2_2 U5376 (.A(net26981), .B(net43702), .Y(n4277));
sg13g2_nand2_2 U5377 (.A(keysched_new_key_o_30), .B(net24849), .Y(n2028));
sg13g2_nand2_2 U5378 (.A(keysched_new_key_o_11), .B(net24857), .Y(n2193));
sg13g2_nor2_2 U5379 (.A(net39214), .B(n4230), .Y(n4280));
sg13g2_nand2_2 U5380 (.A(n4280), .B(n4279), .Y(n4282));
sg13g2_inv_4 U5381 (.A(n3697), .Y(N1123));
sg13g2_nand2_2 U5382 (.A(three_0), .B(net25928), .Y(n3692));
sg13g2_inv_4 U5383 (.A(net26529), .Y(net27467));
sg13g2_xnor2_1 U5384 (.A(keysched_new_key_o_22), .B(addroundkey_data_i_22), .Y(n191));
sg13g2_inv_4 U5385 (.A(N1620), .Y(N1617));
sg13g2_o21ai_1 U5386 (.A1(net24801), .A2(n1034), .B1(n2033), .Y(keysched_last_key_i_26));
sg13g2_inv_4 U5387 (.A(net24881), .Y(net24875));
sg13g2_nand2_2 U5388 (.A(N29), .B(N1610), .Y(n4284));
sg13g2_nand2_2 U5389 (.A(addroundkey_ready_o), .B(decrypt_i), .Y(n3705));
sg13g2_a21oi_2 U5390 (.A1(n4312), .A2(n3397), .B1(n3398), .Y(n3396));
sg13g2_nand2_2 U5391 (.A(keysched_new_key_o_26), .B(net24863), .Y(n2033));
sg13g2_nand2_2 U5392 (.A(n830), .B(n4285), .Y(sbox_data_i_1));
sg13g2_nand2_2 U5393 (.A(keysched_new_key_o_24), .B(net26430), .Y(n2035));
sg13g2_nand2_2 U5394 (.A(n4286), .B(n2109), .Y(keysched_last_key_i_15));
sg13g2_o21ai_1 U5396 (.A1(n4221), .A2(n882), .B1(n1995), .Y(keysched_last_key_i_60));
sg13g2_o21ai_1 U5397 (.A1(net24795), .A2(n1938), .B1(n1939), .Y(keysched_last_key_i_89));
sg13g2_nand2_2 U5398 (.A(data_o_84_), .B(n4320), .Y(n594));
sg13g2_nand2_2 U5399 (.A(n832), .B(n4287), .Y(sbox_data_i_0));
sg13g2_nand2_2 U5400 (.A(keysched_new_key_o_191), .B(net24845), .Y(n2043));
sg13g2_o21ai_1 U5401 (.A1(net26210), .A2(n862), .B1(n1958), .Y(keysched_last_key_i_7));
sg13g2_o21ai_1 U5402 (.A1(n4326), .A2(n639), .B1(n640), .Y(subbytes_data_i_63));
sg13g2_inv_4 U5403 (.A(n4148), .Y(n4149));
sg13g2_nand2_2 U5404 (.A(n818), .B(n4290), .Y(sbox_data_i_7));
sg13g2_inv_4 U5405 (.A(N1593), .Y(N1594));
sg13g2_xnor2_1 U5406 (.A(net25928), .B(addroundkey_round_1), .Y(r371_n17));
sg13g2_o21ai_1 U5407 (.A1(n4221), .A2(n2221), .B1(n2222), .Y(keysched_last_key_i_106));
sg13g2_nand2_2 U5408 (.A(n4252), .B(subbytes_sbox_data_o_4), .Y(n4291));
sg13g2_nand2_2 U5409 (.A(n824), .B(n4291), .Y(sbox_data_i_4));
sg13g2_o21ai_1 U5410 (.A1(n4332), .A2(n3415), .B1(n3416), .Y(addroundkey_data_i_109));
sg13g2_a21oi_2 U5411 (.A1(n4312), .A2(n3417), .B1(n3418), .Y(n3416));
sg13g2_inv_4 U5412 (.A(n560), .Y(n4295));
sg13g2_o21ai_1 U5413 (.A1(n4326), .A2(n637), .B1(n638), .Y(subbytes_data_i_64));
sg13g2_o21ai_1 U5414 (.A1(n4329), .A2(n759), .B1(n760), .Y(subbytes_data_i_124));
sg13g2_nand2_2 U5415 (.A(n4212), .B(N1537), .Y(n1909));
sg13g2_o21ai_1 U5416 (.A1(n4325), .A2(n605), .B1(n606), .Y(subbytes_data_i_79));
sg13g2_nand2_2 U5417 (.A(data_o_47_), .B(n4319), .Y(n676));
sg13g2_a21oi_2 U5418 (.A1(net24687), .A2(N818), .B1(n1472), .Y(n1471));
sg13g2_nor2_2 U5419 (.A(r372_n17), .B(r372_n15), .Y(r372_n13));
sg13g2_nand2_2 U5420 (.A(r372_n13), .B(r372_n19), .Y(r372_n12));
sg13g2_o21ai_1 U5421 (.A1(net24783), .A2(n858), .B1(n1937), .Y(keysched_last_key_i_8));
sg13g2_nand2_2 U5422 (.A(N1323), .B(N1118), .Y(n3725));
sg13g2_o21ai_1 U5423 (.A1(net24795), .A2(n2135), .B1(n2136), .Y(keysched_last_key_i_147));
sg13g2_o21ai_1 U5424 (.A1(n4221), .A2(n2137), .B1(n2138), .Y(keysched_last_key_i_146));
sg13g2_o21ai_1 U5425 (.A1(net24787), .A2(n1058), .B1(n2039), .Y(keysched_last_key_i_20));
sg13g2_nand2_2 U5426 (.A(keysched_sbox_data_o_7), .B(net26029), .Y(n818));
sg13g2_o21ai_1 U5427 (.A1(net26188), .A2(n2229), .B1(n2230), .Y(keysched_last_key_i_102));
sg13g2_o21ai_1 U5428 (.A1(net24795), .A2(n2231), .B1(n2232), .Y(keysched_last_key_i_101));
sg13g2_inv_4 U5429 (.A(net24875), .Y(net24845));
sg13g2_nand2_2 U5430 (.A(keysched_sbox_data_o_3), .B(net26029), .Y(n826));
sg13g2_nand2_2 U5431 (.A(n554), .B(n4166), .Y(n851));
sg13g2_inv_4 U5432 (.A(net44819), .Y(net26864));
sg13g2_nand2_2 U5433 (.A(data_o_64_), .B(n4321), .Y(n638));
sg13g2_nand2_2 U5434 (.A(n4321), .B(data_o_123_), .Y(n762));
sg13g2_o21ai_1 U5435 (.A1(n4325), .A2(n575), .B1(n576), .Y(subbytes_data_i_92));
sg13g2_o21ai_1 U5436 (.A1(n4326), .A2(n675), .B1(n676), .Y(subbytes_data_i_47));
sg13g2_o21ai_1 U5437 (.A1(n4328), .A2(n645), .B1(n646), .Y(subbytes_data_i_60));
sg13g2_nand2_2 U5438 (.A(n4293), .B(mixcol_data_o_75), .Y(n4297));
sg13g2_nand2_2 U5439 (.A(data_o_15_), .B(n4316), .Y(n746));
sg13g2_nand2_2 U5440 (.A(data_o_59_), .B(n4323), .Y(n650));
sg13g2_o21ai_1 U5441 (.A1(n4329), .A2(n629), .B1(n630), .Y(subbytes_data_i_68));
sg13g2_nand2_2 U5442 (.A(data_o_85_), .B(n4319), .Y(n592));
sg13g2_o21ai_1 U5443 (.A1(n4330), .A2(n591), .B1(n592), .Y(subbytes_data_i_85));
sg13g2_nand2_2 U5444 (.A(data_o_76_), .B(n4323), .Y(n612));
sg13g2_nand2_2 U5445 (.A(data_o_92_), .B(n4321), .Y(n576));
sg13g2_o21ai_1 U5446 (.A1(n4325), .A2(n611), .B1(n612), .Y(subbytes_data_i_76));
sg13g2_nand2_2 U5447 (.A(n4299), .B(n2040), .Y(keysched_last_key_i_1));
sg13g2_nand2_2 U5448 (.A(keysched_new_key_o_1), .B(net24863), .Y(n2040));
sg13g2_nand2_2 U5449 (.A(net26529), .B(subbytes_sbox_data_o_3), .Y(n4306));
sg13g2_inv_4 U5450 (.A(n4295), .Y(n4319));
sg13g2_o21ai_1 U5451 (.A1(n4327), .A2(n745), .B1(n746), .Y(subbytes_data_i_15));
sg13g2_o21ai_1 U5452 (.A1(net24795), .A2(n1967), .B1(n1968), .Y(keysched_last_key_i_75));
sg13g2_o21ai_1 U5453 (.A1(net26188), .A2(n2233), .B1(n2234), .Y(keysched_last_key_i_100));
sg13g2_nand2_2 U5454 (.A(keysched_sbox_data_o_1), .B(net26029), .Y(n830));
sg13g2_o21ai_1 U5455 (.A1(n4329), .A2(n585), .B1(n586), .Y(subbytes_data_i_88));
sg13g2_o21ai_1 U5456 (.A1(n4327), .A2(n753), .B1(n754), .Y(subbytes_data_i_127));
sg13g2_o21ai_1 U5457 (.A1(n4327), .A2(n571), .B1(n572), .Y(subbytes_data_i_94));
sg13g2_nand2_2 U5458 (.A(n4304), .B(net44340), .Y(n4301));
sg13g2_nand2_2 U5459 (.A(n4300), .B(n4301), .Y(r371_n10));
sg13g2_nand2_2 U5460 (.A(n4145), .B(N1), .Y(n4302));
sg13g2_nand2_2 U5461 (.A(n4146), .B(net47654), .Y(n4303));
sg13g2_nand2_2 U5462 (.A(n4302), .B(n4303), .Y(n4304));
sg13g2_o21ai_1 U5463 (.A1(n4211), .A2(n2057), .B1(n2058), .Y(keysched_last_key_i_184));
sg13g2_o21ai_1 U5464 (.A1(net24693), .A2(n938), .B1(n939), .Y(next_last_key_half_48));
sg13g2_o21ai_1 U5465 (.A1(net24791), .A2(n1971), .B1(n1972), .Y(keysched_last_key_i_73));
sg13g2_o21ai_1 U5466 (.A1(net24795), .A2(n1990), .B1(n1991), .Y(keysched_last_key_i_64));
sg13g2_a21oi_2 U5467 (.A1(data_i_38_), .A2(n4308), .B1(n2934), .Y(n2933));
sg13g2_o21ai_1 U5468 (.A1(n4328), .A2(n693), .B1(n694), .Y(subbytes_data_i_39));
sg13g2_nand2_2 U5469 (.A(data_o_39_), .B(n4298), .Y(n694));
sg13g2_a21oi_2 U5470 (.A1(n4315), .A2(n3421), .B1(n3422), .Y(n3420));
sg13g2_o21ai_1 U5471 (.A1(n4330), .A2(n3419), .B1(n3423), .Y(n3421));
sg13g2_nand2_2 U5472 (.A(keysched_new_key_o_25), .B(net24863), .Y(n2034));
sg13g2_o21ai_1 U5473 (.A1(n4327), .A2(n767), .B1(n768), .Y(subbytes_data_i_120));
sg13g2_nand2_2 U5474 (.A(n4293), .B(mixcol_data_o_93), .Y(n4305));
sg13g2_nand2_2 U5475 (.A(n574), .B(n4305), .Y(subbytes_data_i_93));
sg13g2_o21ai_1 U5476 (.A1(n4328), .A2(n627), .B1(n628), .Y(subbytes_data_i_69));
sg13g2_o21ai_1 U5477 (.A1(n4325), .A2(n619), .B1(n620), .Y(subbytes_data_i_72));
sg13g2_o21ai_1 U5478 (.A1(net24787), .A2(n1018), .B1(n2029), .Y(keysched_last_key_i_2));
sg13g2_inv_4 U5479 (.A(n4163), .Y(n4321));
sg13g2_inv_4 U5480 (.A(n4324), .Y(n4318));
sg13g2_inv_4 U5481 (.A(n4163), .Y(n4317));
sg13g2_inv_4 U5482 (.A(n4324), .Y(n4316));
sg13g2_o21ai_1 U5483 (.A1(n4325), .A2(n609), .B1(n610), .Y(subbytes_data_i_77));
sg13g2_nand2_2 U5484 (.A(keysched_new_key_o_21), .B(net24847), .Y(n2038));
sg13g2_nand2_2 U5485 (.A(n826), .B(n4306), .Y(sbox_data_i_3));
sg13g2_nand2_2 U5486 (.A(keysched_sbox_data_o_0), .B(net27467), .Y(n832));
sg13g2_nand2_2 U5487 (.A(keysched_new_key_o_13), .B(net24857), .Y(n2151));
sg13g2_o21ai_1 U5488 (.A1(net26188), .A2(n1923), .B1(n1924), .Y(keysched_last_key_i_96));
sg13g2_nand2_2 U5489 (.A(keysched_sbox_data_o_4), .B(net26029), .Y(n824));
sg13g2_inv_4 U5490 (.A(net38935), .Y(net24687));
sg13g2_inv_4 U5491 (.A(net38935), .Y(net24685));
sg13g2_nand2_2 U5492 (.A(n4284), .B(n1904), .Y(n560));
sg13g2_mux2_2 U5493 (.A0(net25972), .A1(next_round_0), .S(N1567), .X(n4129));
sg13g2_nand2_2 U5494 (.A(net25972), .B(n3684), .Y(N1589));
sg13g2_nand2_2 U5495 (.A(net25972), .B(n3676), .Y(N1602));
sg13g2_nand2_2 U5496 (.A(n4162), .B(n4229), .Y(n1904));
sg13g2_mux2_2 U5497 (.A0(net47653), .A1(next_round_3), .S(N1567), .X(n4133));
sg13g2_inv_4 U5498 (.A(n1134), .Y(net24693));
sg13g2_nand2_2 U5499 (.A(net26537), .B(net47654), .Y(N1600));
sg13g2_mux2_2 U5500 (.A0(r371_n27), .A1(next_round_1), .S(N1567), .X(n4130));
sg13g2_a21oi_2 U5501 (.A1(N313), .A2(state), .B1(n1775), .Y(mixcol_start_i));
sg13g2_mux2_2 U5502 (.A0(net26538), .A1(next_round_2), .S(N1567), .X(n4131));
sg13g2_nand2_2 U5503 (.A(n4160), .B(n4157), .Y(n1905));
sg13g2_xnor2_1 U5504 (.A(keysched_new_key_o_100), .B(addroundkey_data_i_100), .Y(n269));
sg13g2_xnor2_1 U5505 (.A(keysched_new_key_o_101), .B(addroundkey_data_i_101), .Y(n270));
sg13g2_xnor2_1 U5506 (.A(keysched_new_key_o_102), .B(addroundkey_data_i_102), .Y(n271));
sg13g2_inv_4 U5507 (.A(net38935), .Y(net24689));
sg13g2_xnor2_1 U5508 (.A(keysched_new_key_o_103), .B(addroundkey_data_i_103), .Y(n272));
sg13g2_xnor2_1 U5509 (.A(keysched_new_key_o_104), .B(addroundkey_data_i_104), .Y(n273));
sg13g2_xnor2_1 U5510 (.A(keysched_new_key_o_105), .B(addroundkey_data_i_105), .Y(n274));
sg13g2_xnor2_1 U5511 (.A(keysched_new_key_o_106), .B(addroundkey_data_i_106), .Y(n275));
sg13g2_xnor2_1 U5512 (.A(keysched_new_key_o_107), .B(addroundkey_data_i_107), .Y(n276));
sg13g2_xnor2_1 U5513 (.A(keysched_new_key_o_108), .B(addroundkey_data_i_108), .Y(n277));
sg13g2_xnor2_1 U5514 (.A(keysched_new_key_o_109), .B(addroundkey_data_i_109), .Y(n278));
sg13g2_xnor2_1 U5515 (.A(keysched_new_key_o_10), .B(addroundkey_data_i_10), .Y(n179));
sg13g2_xnor2_1 U5516 (.A(keysched_new_key_o_110), .B(addroundkey_data_i_110), .Y(n279));
sg13g2_xnor2_1 U5517 (.A(keysched_new_key_o_111), .B(addroundkey_data_i_111), .Y(n280));
sg13g2_xnor2_1 U5518 (.A(keysched_new_key_o_112), .B(addroundkey_data_i_112), .Y(n281));
sg13g2_xnor2_1 U5519 (.A(keysched_new_key_o_113), .B(addroundkey_data_i_113), .Y(n282));
sg13g2_xnor2_1 U5520 (.A(keysched_new_key_o_114), .B(addroundkey_data_i_114), .Y(n283));
sg13g2_xnor2_1 U5521 (.A(keysched_new_key_o_115), .B(addroundkey_data_i_115), .Y(n284));
sg13g2_xnor2_1 U5522 (.A(keysched_new_key_o_116), .B(addroundkey_data_i_116), .Y(n285));
sg13g2_xnor2_1 U5523 (.A(keysched_new_key_o_117), .B(addroundkey_data_i_117), .Y(n286));
sg13g2_xnor2_1 U5524 (.A(keysched_new_key_o_118), .B(addroundkey_data_i_118), .Y(n287));
sg13g2_xnor2_1 U5525 (.A(keysched_new_key_o_119), .B(addroundkey_data_i_119), .Y(n288));
sg13g2_xnor2_1 U5526 (.A(keysched_new_key_o_11), .B(addroundkey_data_i_11), .Y(n180));
sg13g2_xnor2_1 U5527 (.A(keysched_new_key_o_120), .B(addroundkey_data_i_120), .Y(n289));
sg13g2_xnor2_1 U5528 (.A(keysched_new_key_o_121), .B(addroundkey_data_i_121), .Y(n290));
sg13g2_xnor2_1 U5529 (.A(keysched_new_key_o_122), .B(addroundkey_data_i_122), .Y(n291));
sg13g2_xnor2_1 U5530 (.A(keysched_new_key_o_123), .B(addroundkey_data_i_123), .Y(n292));
sg13g2_xnor2_1 U5531 (.A(keysched_new_key_o_124), .B(addroundkey_data_i_124), .Y(n293));
sg13g2_xnor2_1 U5532 (.A(keysched_new_key_o_125), .B(addroundkey_data_i_125), .Y(n294));
sg13g2_xnor2_1 U5533 (.A(keysched_new_key_o_126), .B(addroundkey_data_i_126), .Y(n295));
sg13g2_xnor2_1 U5534 (.A(keysched_new_key_o_127), .B(addroundkey_data_i_127), .Y(n296));
sg13g2_xnor2_1 U5535 (.A(keysched_new_key_o_12), .B(addroundkey_data_i_12), .Y(n181));
sg13g2_xnor2_1 U5536 (.A(keysched_new_key_o_13), .B(addroundkey_data_i_13), .Y(n182));
sg13g2_xnor2_1 U5537 (.A(keysched_new_key_o_14), .B(addroundkey_data_i_14), .Y(n183));
sg13g2_xnor2_1 U5538 (.A(keysched_new_key_o_15), .B(addroundkey_data_i_15), .Y(n184));
sg13g2_xnor2_1 U5539 (.A(keysched_new_key_o_16), .B(addroundkey_data_i_16), .Y(n185));
sg13g2_xnor2_1 U5540 (.A(keysched_new_key_o_17), .B(addroundkey_data_i_17), .Y(n186));
sg13g2_xnor2_1 U5541 (.A(keysched_new_key_o_18), .B(addroundkey_data_i_18), .Y(n187));
sg13g2_xnor2_1 U5542 (.A(keysched_new_key_o_19), .B(addroundkey_data_i_19), .Y(n188));
sg13g2_xnor2_1 U5543 (.A(keysched_new_key_o_1), .B(addroundkey_data_i_1), .Y(n170));
sg13g2_xnor2_1 U5544 (.A(keysched_new_key_o_20), .B(addroundkey_data_i_20), .Y(n189));
sg13g2_xnor2_1 U5545 (.A(keysched_new_key_o_21), .B(addroundkey_data_i_21), .Y(n190));
sg13g2_xnor2_1 U5546 (.A(keysched_new_key_o_23), .B(addroundkey_data_i_23), .Y(n192));
sg13g2_xnor2_1 U5547 (.A(keysched_new_key_o_24), .B(addroundkey_data_i_24), .Y(n193));
sg13g2_xnor2_1 U5548 (.A(keysched_new_key_o_25), .B(addroundkey_data_i_25), .Y(n194));
sg13g2_xnor2_1 U5549 (.A(keysched_new_key_o_26), .B(addroundkey_data_i_26), .Y(n195));
sg13g2_xnor2_1 U5550 (.A(keysched_new_key_o_27), .B(addroundkey_data_i_27), .Y(n196));
sg13g2_xnor2_1 U5551 (.A(keysched_new_key_o_28), .B(addroundkey_data_i_28), .Y(n197));
sg13g2_xnor2_1 U5552 (.A(keysched_new_key_o_29), .B(addroundkey_data_i_29), .Y(n198));
sg13g2_xnor2_1 U5553 (.A(keysched_new_key_o_2), .B(addroundkey_data_i_2), .Y(n171));
sg13g2_xnor2_1 U5554 (.A(keysched_new_key_o_30), .B(addroundkey_data_i_30), .Y(n199));
sg13g2_xnor2_1 U5555 (.A(keysched_new_key_o_31), .B(addroundkey_data_i_31), .Y(n200));
sg13g2_xnor2_1 U5556 (.A(keysched_new_key_o_32), .B(addroundkey_data_i_32), .Y(n201));
sg13g2_xnor2_1 U5557 (.A(keysched_new_key_o_33), .B(addroundkey_data_i_33), .Y(n202));
sg13g2_xnor2_1 U5558 (.A(keysched_new_key_o_34), .B(addroundkey_data_i_34), .Y(n203));
sg13g2_xnor2_1 U5559 (.A(keysched_new_key_o_35), .B(addroundkey_data_i_35), .Y(n204));
sg13g2_xnor2_1 U5560 (.A(keysched_new_key_o_36), .B(addroundkey_data_i_36), .Y(n205));
sg13g2_xnor2_1 U5561 (.A(keysched_new_key_o_37), .B(addroundkey_data_i_37), .Y(n206));
sg13g2_xnor2_1 U5562 (.A(keysched_new_key_o_38), .B(addroundkey_data_i_38), .Y(n207));
sg13g2_xnor2_1 U5563 (.A(keysched_new_key_o_39), .B(addroundkey_data_i_39), .Y(n208));
sg13g2_xnor2_1 U5564 (.A(keysched_new_key_o_3), .B(addroundkey_data_i_3), .Y(n172));
sg13g2_xnor2_1 U5565 (.A(keysched_new_key_o_40), .B(addroundkey_data_i_40), .Y(n209));
sg13g2_xnor2_1 U5566 (.A(keysched_new_key_o_41), .B(addroundkey_data_i_41), .Y(n210));
sg13g2_xnor2_1 U5567 (.A(keysched_new_key_o_42), .B(addroundkey_data_i_42), .Y(n211));
sg13g2_xnor2_1 U5568 (.A(keysched_new_key_o_43), .B(addroundkey_data_i_43), .Y(n212));
sg13g2_xnor2_1 U5569 (.A(keysched_new_key_o_44), .B(addroundkey_data_i_44), .Y(n213));
sg13g2_xnor2_1 U5570 (.A(keysched_new_key_o_45), .B(addroundkey_data_i_45), .Y(n214));
sg13g2_xnor2_1 U5571 (.A(keysched_new_key_o_46), .B(addroundkey_data_i_46), .Y(n215));
sg13g2_xnor2_1 U5572 (.A(keysched_new_key_o_47), .B(addroundkey_data_i_47), .Y(n216));
sg13g2_xnor2_1 U5573 (.A(keysched_new_key_o_48), .B(addroundkey_data_i_48), .Y(n217));
sg13g2_xnor2_1 U5574 (.A(keysched_new_key_o_49), .B(addroundkey_data_i_49), .Y(n218));
sg13g2_xnor2_1 U5575 (.A(keysched_new_key_o_4), .B(addroundkey_data_i_4), .Y(n173));
sg13g2_xnor2_1 U5576 (.A(keysched_new_key_o_50), .B(addroundkey_data_i_50), .Y(n219));
sg13g2_xnor2_1 U5577 (.A(keysched_new_key_o_51), .B(addroundkey_data_i_51), .Y(n220));
sg13g2_xnor2_1 U5578 (.A(keysched_new_key_o_52), .B(addroundkey_data_i_52), .Y(n221));
sg13g2_xnor2_1 U5579 (.A(keysched_new_key_o_53), .B(addroundkey_data_i_53), .Y(n222));
sg13g2_xnor2_1 U5580 (.A(keysched_new_key_o_54), .B(addroundkey_data_i_54), .Y(n223));
sg13g2_xnor2_1 U5581 (.A(keysched_new_key_o_55), .B(addroundkey_data_i_55), .Y(n224));
sg13g2_xnor2_1 U5582 (.A(keysched_new_key_o_56), .B(addroundkey_data_i_56), .Y(n225));
sg13g2_xnor2_1 U5583 (.A(keysched_new_key_o_57), .B(addroundkey_data_i_57), .Y(n226));
sg13g2_xnor2_1 U5584 (.A(keysched_new_key_o_58), .B(addroundkey_data_i_58), .Y(n227));
sg13g2_xnor2_1 U5585 (.A(keysched_new_key_o_59), .B(addroundkey_data_i_59), .Y(n228));
sg13g2_xnor2_1 U5586 (.A(keysched_new_key_o_5), .B(addroundkey_data_i_5), .Y(n174));
sg13g2_xnor2_1 U5587 (.A(keysched_new_key_o_60), .B(addroundkey_data_i_60), .Y(n229));
sg13g2_xnor2_1 U5588 (.A(keysched_new_key_o_61), .B(addroundkey_data_i_61), .Y(n230));
sg13g2_xnor2_1 U5589 (.A(keysched_new_key_o_62), .B(addroundkey_data_i_62), .Y(n231));
sg13g2_xnor2_1 U5590 (.A(keysched_new_key_o_63), .B(addroundkey_data_i_63), .Y(n232));
sg13g2_xnor2_1 U5591 (.A(keysched_new_key_o_64), .B(addroundkey_data_i_64), .Y(n233));
sg13g2_xnor2_1 U5592 (.A(keysched_new_key_o_65), .B(addroundkey_data_i_65), .Y(n234));
sg13g2_xnor2_1 U5593 (.A(keysched_new_key_o_66), .B(addroundkey_data_i_66), .Y(n235));
sg13g2_xnor2_1 U5594 (.A(keysched_new_key_o_67), .B(addroundkey_data_i_67), .Y(n236));
sg13g2_xnor2_1 U5595 (.A(keysched_new_key_o_68), .B(addroundkey_data_i_68), .Y(n237));
sg13g2_xnor2_1 U5596 (.A(keysched_new_key_o_69), .B(addroundkey_data_i_69), .Y(n238));
sg13g2_xnor2_1 U5597 (.A(keysched_new_key_o_6), .B(addroundkey_data_i_6), .Y(n175));
sg13g2_xnor2_1 U5598 (.A(keysched_new_key_o_70), .B(addroundkey_data_i_70), .Y(n239));
sg13g2_xnor2_1 U5599 (.A(keysched_new_key_o_71), .B(addroundkey_data_i_71), .Y(n240));
sg13g2_xnor2_1 U5600 (.A(keysched_new_key_o_72), .B(addroundkey_data_i_72), .Y(n241));
sg13g2_xnor2_1 U5601 (.A(keysched_new_key_o_74), .B(addroundkey_data_i_74), .Y(n243));
sg13g2_xnor2_1 U5602 (.A(keysched_new_key_o_75), .B(addroundkey_data_i_75), .Y(n244));
sg13g2_xnor2_1 U5603 (.A(keysched_new_key_o_76), .B(addroundkey_data_i_76), .Y(n245));
sg13g2_xnor2_1 U5604 (.A(keysched_new_key_o_77), .B(addroundkey_data_i_77), .Y(n246));
sg13g2_xnor2_1 U5605 (.A(keysched_new_key_o_78), .B(addroundkey_data_i_78), .Y(n247));
sg13g2_xnor2_1 U5606 (.A(keysched_new_key_o_79), .B(addroundkey_data_i_79), .Y(n248));
sg13g2_xnor2_1 U5607 (.A(keysched_new_key_o_7), .B(addroundkey_data_i_7), .Y(n176));
sg13g2_xnor2_1 U5608 (.A(keysched_new_key_o_80), .B(addroundkey_data_i_80), .Y(n249));
sg13g2_xnor2_1 U5609 (.A(keysched_new_key_o_81), .B(addroundkey_data_i_81), .Y(n250));
sg13g2_xnor2_1 U5610 (.A(keysched_new_key_o_82), .B(addroundkey_data_i_82), .Y(n251));
sg13g2_xnor2_1 U5611 (.A(keysched_new_key_o_83), .B(addroundkey_data_i_83), .Y(n252));
sg13g2_xnor2_1 U5612 (.A(keysched_new_key_o_84), .B(addroundkey_data_i_84), .Y(n253));
sg13g2_xnor2_1 U5613 (.A(keysched_new_key_o_85), .B(addroundkey_data_i_85), .Y(n254));
sg13g2_xnor2_1 U5614 (.A(keysched_new_key_o_86), .B(addroundkey_data_i_86), .Y(n255));
sg13g2_xnor2_1 U5615 (.A(keysched_new_key_o_87), .B(addroundkey_data_i_87), .Y(n256));
sg13g2_xnor2_1 U5616 (.A(keysched_new_key_o_88), .B(addroundkey_data_i_88), .Y(n257));
sg13g2_xnor2_1 U5617 (.A(keysched_new_key_o_89), .B(addroundkey_data_i_89), .Y(n258));
sg13g2_xnor2_1 U5618 (.A(keysched_new_key_o_8), .B(addroundkey_data_i_8), .Y(n177));
sg13g2_xnor2_1 U5619 (.A(keysched_new_key_o_90), .B(addroundkey_data_i_90), .Y(n259));
sg13g2_xnor2_1 U5620 (.A(keysched_new_key_o_91), .B(addroundkey_data_i_91), .Y(n260));
sg13g2_xnor2_1 U5621 (.A(keysched_new_key_o_92), .B(addroundkey_data_i_92), .Y(n261));
sg13g2_xnor2_1 U5622 (.A(keysched_new_key_o_93), .B(addroundkey_data_i_93), .Y(n262));
sg13g2_xnor2_1 U5623 (.A(keysched_new_key_o_94), .B(addroundkey_data_i_94), .Y(n263));
sg13g2_xnor2_1 U5624 (.A(keysched_new_key_o_95), .B(addroundkey_data_i_95), .Y(n264));
sg13g2_xnor2_1 U5625 (.A(keysched_new_key_o_96), .B(addroundkey_data_i_96), .Y(n265));
sg13g2_xnor2_1 U5626 (.A(keysched_new_key_o_97), .B(addroundkey_data_i_97), .Y(n266));
sg13g2_xnor2_1 U5627 (.A(keysched_new_key_o_98), .B(addroundkey_data_i_98), .Y(n267));
sg13g2_xnor2_1 U5628 (.A(keysched_new_key_o_99), .B(addroundkey_data_i_99), .Y(n268));
sg13g2_xnor2_1 U5629 (.A(keysched_new_key_o_9), .B(addroundkey_data_i_9), .Y(n178));
sg13g2_xnor2_1 U5630 (.A(keysched_new_key_o_0), .B(addroundkey_data_i_0), .Y(n169));
sg13g2_xnor2_1 U5631 (.A(keysched_new_key_o_73), .B(addroundkey_data_i_73), .Y(n242));
sg13g2_inv_4 U5632 (.A(n3699), .Y(N1121));
sg13g2_inv_4 U5633 (.A(n525), .Y(N757));
sg13g2_xnor2_1 U5634 (.A(key_i_164_), .B(addroundkey_data_i_100), .Y(n525));
sg13g2_inv_4 U5635 (.A(n269), .Y(N1013));
sg13g2_xnor2_1 U5636 (.A(N1378), .B(addroundkey_data_i_100), .Y(n137));
sg13g2_inv_4 U5637 (.A(n526), .Y(N756));
sg13g2_xnor2_1 U5638 (.A(key_i_165_), .B(addroundkey_data_i_101), .Y(n526));
sg13g2_inv_4 U5639 (.A(n270), .Y(N1012));
sg13g2_xnor2_1 U5640 (.A(N1379), .B(addroundkey_data_i_101), .Y(n138));
sg13g2_inv_4 U5641 (.A(n527), .Y(N755));
sg13g2_xnor2_1 U5642 (.A(key_i_166_), .B(addroundkey_data_i_102), .Y(n527));
sg13g2_inv_4 U5643 (.A(n271), .Y(N1011));
sg13g2_xnor2_1 U5644 (.A(N1380), .B(addroundkey_data_i_102), .Y(n139));
sg13g2_inv_4 U5645 (.A(n528), .Y(N754));
sg13g2_xnor2_1 U5646 (.A(key_i_167_), .B(addroundkey_data_i_103), .Y(n528));
sg13g2_inv_4 U5647 (.A(n272), .Y(N1010));
sg13g2_xnor2_1 U5648 (.A(N1381), .B(addroundkey_data_i_103), .Y(n140));
sg13g2_inv_4 U5649 (.A(n273), .Y(N1009));
sg13g2_xnor2_1 U5650 (.A(N1382), .B(addroundkey_data_i_104), .Y(n141));
sg13g2_inv_4 U5651 (.A(n274), .Y(N1008));
sg13g2_xnor2_1 U5652 (.A(N1383), .B(addroundkey_data_i_105), .Y(n142));
sg13g2_inv_4 U5653 (.A(n275), .Y(N1007));
sg13g2_xnor2_1 U5654 (.A(N1384), .B(addroundkey_data_i_106), .Y(n143));
sg13g2_inv_4 U5655 (.A(n276), .Y(N1006));
sg13g2_xnor2_1 U5656 (.A(N1385), .B(addroundkey_data_i_107), .Y(n144));
sg13g2_inv_4 U5657 (.A(n277), .Y(N1005));
sg13g2_xnor2_1 U5658 (.A(N1386), .B(addroundkey_data_i_108), .Y(n145));
sg13g2_inv_4 U5659 (.A(n278), .Y(N1004));
sg13g2_xnor2_1 U5660 (.A(N1387), .B(addroundkey_data_i_109), .Y(n146));
sg13g2_inv_4 U5661 (.A(n179), .Y(N1103));
sg13g2_xnor2_1 U5662 (.A(keysched_new_key_o_138), .B(addroundkey_data_i_10), .Y(n47));
sg13g2_inv_4 U5663 (.A(n279), .Y(N1003));
sg13g2_xnor2_1 U5664 (.A(N1388), .B(addroundkey_data_i_110), .Y(n147));
sg13g2_inv_4 U5665 (.A(n280), .Y(N1002));
sg13g2_xnor2_1 U5666 (.A(N1389), .B(addroundkey_data_i_111), .Y(n148));
sg13g2_inv_4 U5667 (.A(n281), .Y(N1001));
sg13g2_xnor2_1 U5668 (.A(N1390), .B(addroundkey_data_i_112), .Y(n149));
sg13g2_inv_4 U5669 (.A(n282), .Y(N1000));
sg13g2_xnor2_1 U5670 (.A(N1391), .B(addroundkey_data_i_113), .Y(n150));
sg13g2_inv_4 U5671 (.A(n283), .Y(N999));
sg13g2_xnor2_1 U5672 (.A(N1392), .B(addroundkey_data_i_114), .Y(n151));
sg13g2_inv_4 U5673 (.A(n284), .Y(N998));
sg13g2_xnor2_1 U5674 (.A(N1393), .B(addroundkey_data_i_115), .Y(n152));
sg13g2_inv_4 U5675 (.A(n285), .Y(N997));
sg13g2_xnor2_1 U5676 (.A(N1394), .B(addroundkey_data_i_116), .Y(n153));
sg13g2_inv_4 U5677 (.A(n286), .Y(N996));
sg13g2_xnor2_1 U5678 (.A(N1395), .B(addroundkey_data_i_117), .Y(n154));
sg13g2_inv_4 U5679 (.A(n287), .Y(N995));
sg13g2_xnor2_1 U5680 (.A(N1396), .B(addroundkey_data_i_118), .Y(n155));
sg13g2_inv_4 U5681 (.A(n288), .Y(N994));
sg13g2_xnor2_1 U5682 (.A(N1397), .B(addroundkey_data_i_119), .Y(n156));
sg13g2_inv_4 U5683 (.A(n180), .Y(N1102));
sg13g2_xnor2_1 U5684 (.A(keysched_new_key_o_139), .B(addroundkey_data_i_11), .Y(n48));
sg13g2_inv_4 U5685 (.A(n289), .Y(N993));
sg13g2_xnor2_1 U5686 (.A(N1398), .B(addroundkey_data_i_120), .Y(n157));
sg13g2_inv_4 U5687 (.A(n290), .Y(N992));
sg13g2_xnor2_1 U5688 (.A(N1399), .B(addroundkey_data_i_121), .Y(n158));
sg13g2_inv_4 U5689 (.A(n291), .Y(N991));
sg13g2_xnor2_1 U5690 (.A(N1400), .B(addroundkey_data_i_122), .Y(n159));
sg13g2_inv_4 U5691 (.A(n292), .Y(N990));
sg13g2_xnor2_1 U5692 (.A(N1401), .B(addroundkey_data_i_123), .Y(n160));
sg13g2_inv_4 U5693 (.A(n549), .Y(N733));
sg13g2_xnor2_1 U5694 (.A(key_i_188_), .B(addroundkey_data_i_124), .Y(n549));
sg13g2_inv_4 U5695 (.A(n293), .Y(N989));
sg13g2_xnor2_1 U5696 (.A(N1402), .B(addroundkey_data_i_124), .Y(n161));
sg13g2_inv_4 U5697 (.A(n550), .Y(N732));
sg13g2_xnor2_1 U5698 (.A(key_i_189_), .B(addroundkey_data_i_125), .Y(n550));
sg13g2_inv_4 U5699 (.A(n294), .Y(N988));
sg13g2_xnor2_1 U5700 (.A(N1403), .B(addroundkey_data_i_125), .Y(n162));
sg13g2_inv_4 U5701 (.A(n551), .Y(N731));
sg13g2_xnor2_1 U5702 (.A(key_i_190_), .B(addroundkey_data_i_126), .Y(n551));
sg13g2_inv_4 U5703 (.A(n295), .Y(N987));
sg13g2_xnor2_1 U5704 (.A(N1404), .B(addroundkey_data_i_126), .Y(n163));
sg13g2_inv_4 U5705 (.A(n552), .Y(N730));
sg13g2_xnor2_1 U5706 (.A(key_i_191_), .B(addroundkey_data_i_127), .Y(n552));
sg13g2_inv_4 U5707 (.A(n296), .Y(N986));
sg13g2_xnor2_1 U5708 (.A(N1405), .B(addroundkey_data_i_127), .Y(n164));
sg13g2_inv_4 U5709 (.A(n437), .Y(N845));
sg13g2_xnor2_1 U5710 (.A(key_i_76_), .B(addroundkey_data_i_12), .Y(n437));
sg13g2_inv_4 U5711 (.A(n181), .Y(N1101));
sg13g2_xnor2_1 U5712 (.A(keysched_new_key_o_140), .B(addroundkey_data_i_12), .Y(n49));
sg13g2_inv_4 U5713 (.A(n438), .Y(N844));
sg13g2_xnor2_1 U5714 (.A(key_i_77_), .B(addroundkey_data_i_13), .Y(n438));
sg13g2_inv_4 U5715 (.A(n182), .Y(N1100));
sg13g2_xnor2_1 U5716 (.A(keysched_new_key_o_141), .B(addroundkey_data_i_13), .Y(n50));
sg13g2_inv_4 U5717 (.A(n439), .Y(N843));
sg13g2_xnor2_1 U5718 (.A(key_i_78_), .B(addroundkey_data_i_14), .Y(n439));
sg13g2_inv_4 U5719 (.A(n183), .Y(N1099));
sg13g2_xnor2_1 U5720 (.A(keysched_new_key_o_142), .B(addroundkey_data_i_14), .Y(n51));
sg13g2_inv_4 U5721 (.A(n440), .Y(N842));
sg13g2_xnor2_1 U5722 (.A(key_i_79_), .B(addroundkey_data_i_15), .Y(n440));
sg13g2_inv_4 U5723 (.A(n184), .Y(N1098));
sg13g2_xnor2_1 U5724 (.A(keysched_new_key_o_143), .B(addroundkey_data_i_15), .Y(n52));
sg13g2_inv_4 U5725 (.A(n441), .Y(N841));
sg13g2_xnor2_1 U5726 (.A(key_i_80_), .B(addroundkey_data_i_16), .Y(n441));
sg13g2_inv_4 U5727 (.A(n185), .Y(N1097));
sg13g2_xnor2_1 U5728 (.A(keysched_new_key_o_144), .B(addroundkey_data_i_16), .Y(n53));
sg13g2_inv_4 U5729 (.A(n442), .Y(N840));
sg13g2_xnor2_1 U5730 (.A(key_i_81_), .B(addroundkey_data_i_17), .Y(n442));
sg13g2_inv_4 U5731 (.A(n186), .Y(N1096));
sg13g2_xnor2_1 U5732 (.A(keysched_new_key_o_145), .B(addroundkey_data_i_17), .Y(n54));
sg13g2_inv_4 U5733 (.A(n443), .Y(N839));
sg13g2_xnor2_1 U5734 (.A(key_i_82_), .B(addroundkey_data_i_18), .Y(n443));
sg13g2_inv_4 U5735 (.A(n187), .Y(N1095));
sg13g2_xnor2_1 U5736 (.A(keysched_new_key_o_146), .B(addroundkey_data_i_18), .Y(n55));
sg13g2_inv_4 U5737 (.A(n444), .Y(N838));
sg13g2_xnor2_1 U5738 (.A(key_i_83_), .B(addroundkey_data_i_19), .Y(n444));
sg13g2_inv_4 U5739 (.A(n188), .Y(N1094));
sg13g2_xnor2_1 U5740 (.A(keysched_new_key_o_147), .B(addroundkey_data_i_19), .Y(n56));
sg13g2_inv_4 U5741 (.A(n426), .Y(N856));
sg13g2_xnor2_1 U5742 (.A(key_i_65_), .B(addroundkey_data_i_1), .Y(n426));
sg13g2_inv_4 U5743 (.A(n170), .Y(N1112));
sg13g2_xnor2_1 U5744 (.A(keysched_new_key_o_129), .B(addroundkey_data_i_1), .Y(n38));
sg13g2_inv_4 U5745 (.A(n445), .Y(N837));
sg13g2_xnor2_1 U5746 (.A(key_i_84_), .B(addroundkey_data_i_20), .Y(n445));
sg13g2_inv_4 U5747 (.A(n189), .Y(N1093));
sg13g2_xnor2_1 U5748 (.A(keysched_new_key_o_148), .B(addroundkey_data_i_20), .Y(n57));
sg13g2_inv_4 U5749 (.A(n446), .Y(N836));
sg13g2_xnor2_1 U5750 (.A(key_i_85_), .B(addroundkey_data_i_21), .Y(n446));
sg13g2_inv_4 U5751 (.A(n190), .Y(N1092));
sg13g2_xnor2_1 U5752 (.A(keysched_new_key_o_149), .B(addroundkey_data_i_21), .Y(n58));
sg13g2_inv_4 U5753 (.A(n447), .Y(N835));
sg13g2_xnor2_1 U5754 (.A(key_i_86_), .B(addroundkey_data_i_22), .Y(n447));
sg13g2_inv_4 U5755 (.A(n191), .Y(N1091));
sg13g2_xnor2_1 U5756 (.A(keysched_new_key_o_150), .B(addroundkey_data_i_22), .Y(n59));
sg13g2_inv_4 U5757 (.A(n448), .Y(N834));
sg13g2_xnor2_1 U5758 (.A(key_i_87_), .B(addroundkey_data_i_23), .Y(n448));
sg13g2_inv_4 U5759 (.A(n192), .Y(N1090));
sg13g2_xnor2_1 U5760 (.A(keysched_new_key_o_151), .B(addroundkey_data_i_23), .Y(n60));
sg13g2_inv_4 U5761 (.A(n449), .Y(N833));
sg13g2_xnor2_1 U5762 (.A(key_i_88_), .B(addroundkey_data_i_24), .Y(n449));
sg13g2_inv_4 U5763 (.A(n193), .Y(N1089));
sg13g2_xnor2_1 U5764 (.A(keysched_new_key_o_152), .B(addroundkey_data_i_24), .Y(n61));
sg13g2_inv_4 U5765 (.A(n450), .Y(N832));
sg13g2_xnor2_1 U5766 (.A(key_i_89_), .B(addroundkey_data_i_25), .Y(n450));
sg13g2_inv_4 U5767 (.A(n194), .Y(N1088));
sg13g2_xnor2_1 U5768 (.A(keysched_new_key_o_153), .B(addroundkey_data_i_25), .Y(n62));
sg13g2_inv_4 U5769 (.A(n451), .Y(N831));
sg13g2_xnor2_1 U5770 (.A(key_i_90_), .B(addroundkey_data_i_26), .Y(n451));
sg13g2_inv_4 U5771 (.A(n195), .Y(N1087));
sg13g2_xnor2_1 U5772 (.A(keysched_new_key_o_154), .B(addroundkey_data_i_26), .Y(n63));
sg13g2_inv_4 U5773 (.A(n452), .Y(N830));
sg13g2_xnor2_1 U5774 (.A(key_i_91_), .B(addroundkey_data_i_27), .Y(n452));
sg13g2_inv_4 U5775 (.A(n196), .Y(N1086));
sg13g2_xnor2_1 U5776 (.A(keysched_new_key_o_155), .B(addroundkey_data_i_27), .Y(n64));
sg13g2_inv_4 U5777 (.A(n453), .Y(N829));
sg13g2_xnor2_1 U5778 (.A(key_i_92_), .B(addroundkey_data_i_28), .Y(n453));
sg13g2_inv_4 U5779 (.A(n197), .Y(N1085));
sg13g2_xnor2_1 U5780 (.A(keysched_new_key_o_156), .B(addroundkey_data_i_28), .Y(n65));
sg13g2_inv_4 U5781 (.A(n454), .Y(N828));
sg13g2_xnor2_1 U5782 (.A(key_i_93_), .B(addroundkey_data_i_29), .Y(n454));
sg13g2_inv_4 U5783 (.A(n198), .Y(N1084));
sg13g2_xnor2_1 U5784 (.A(keysched_new_key_o_157), .B(addroundkey_data_i_29), .Y(n66));
sg13g2_inv_4 U5785 (.A(n427), .Y(N855));
sg13g2_xnor2_1 U5786 (.A(key_i_66_), .B(addroundkey_data_i_2), .Y(n427));
sg13g2_inv_4 U5787 (.A(n171), .Y(N1111));
sg13g2_xnor2_1 U5788 (.A(keysched_new_key_o_130), .B(addroundkey_data_i_2), .Y(n39));
sg13g2_inv_4 U5789 (.A(n455), .Y(N827));
sg13g2_xnor2_1 U5790 (.A(key_i_94_), .B(addroundkey_data_i_30), .Y(n455));
sg13g2_inv_4 U5791 (.A(n199), .Y(N1083));
sg13g2_xnor2_1 U5792 (.A(keysched_new_key_o_158), .B(addroundkey_data_i_30), .Y(n67));
sg13g2_inv_4 U5793 (.A(n456), .Y(N826));
sg13g2_xnor2_1 U5794 (.A(key_i_95_), .B(addroundkey_data_i_31), .Y(n456));
sg13g2_inv_4 U5795 (.A(n200), .Y(N1082));
sg13g2_xnor2_1 U5796 (.A(keysched_new_key_o_159), .B(addroundkey_data_i_31), .Y(n68));
sg13g2_inv_4 U5797 (.A(n457), .Y(N825));
sg13g2_xnor2_1 U5798 (.A(key_i_96_), .B(addroundkey_data_i_32), .Y(n457));
sg13g2_inv_4 U5799 (.A(n201), .Y(N1081));
sg13g2_xnor2_1 U5800 (.A(keysched_new_key_o_160), .B(addroundkey_data_i_32), .Y(n69));
sg13g2_inv_4 U5801 (.A(n458), .Y(N824));
sg13g2_xnor2_1 U5802 (.A(key_i_97_), .B(addroundkey_data_i_33), .Y(n458));
sg13g2_inv_4 U5803 (.A(n202), .Y(N1080));
sg13g2_xnor2_1 U5804 (.A(keysched_new_key_o_161), .B(addroundkey_data_i_33), .Y(n70));
sg13g2_inv_4 U5805 (.A(n459), .Y(N823));
sg13g2_xnor2_1 U5806 (.A(key_i_98_), .B(addroundkey_data_i_34), .Y(n459));
sg13g2_inv_4 U5807 (.A(n203), .Y(N1079));
sg13g2_xnor2_1 U5808 (.A(keysched_new_key_o_162), .B(addroundkey_data_i_34), .Y(n71));
sg13g2_inv_4 U5809 (.A(n460), .Y(N822));
sg13g2_xnor2_1 U5810 (.A(key_i_99_), .B(addroundkey_data_i_35), .Y(n460));
sg13g2_inv_4 U5811 (.A(n204), .Y(N1078));
sg13g2_xnor2_1 U5812 (.A(keysched_new_key_o_163), .B(addroundkey_data_i_35), .Y(n72));
sg13g2_inv_4 U5813 (.A(n461), .Y(N821));
sg13g2_xnor2_1 U5814 (.A(key_i_100_), .B(addroundkey_data_i_36), .Y(n461));
sg13g2_inv_4 U5815 (.A(n205), .Y(N1077));
sg13g2_xnor2_1 U5816 (.A(keysched_new_key_o_164), .B(addroundkey_data_i_36), .Y(n73));
sg13g2_inv_4 U5817 (.A(n462), .Y(N820));
sg13g2_xnor2_1 U5818 (.A(key_i_101_), .B(addroundkey_data_i_37), .Y(n462));
sg13g2_inv_4 U5819 (.A(n206), .Y(N1076));
sg13g2_xnor2_1 U5820 (.A(keysched_new_key_o_165), .B(addroundkey_data_i_37), .Y(n74));
sg13g2_inv_4 U5821 (.A(n463), .Y(N819));
sg13g2_xnor2_1 U5822 (.A(key_i_102_), .B(addroundkey_data_i_38), .Y(n463));
sg13g2_inv_4 U5823 (.A(n207), .Y(N1075));
sg13g2_xnor2_1 U5824 (.A(keysched_new_key_o_166), .B(addroundkey_data_i_38), .Y(n75));
sg13g2_inv_4 U5825 (.A(n464), .Y(N818));
sg13g2_xnor2_1 U5826 (.A(key_i_103_), .B(addroundkey_data_i_39), .Y(n464));
sg13g2_inv_4 U5827 (.A(n208), .Y(N1074));
sg13g2_xnor2_1 U5828 (.A(keysched_new_key_o_167), .B(addroundkey_data_i_39), .Y(n76));
sg13g2_inv_4 U5829 (.A(n428), .Y(N854));
sg13g2_xnor2_1 U5830 (.A(key_i_67_), .B(addroundkey_data_i_3), .Y(n428));
sg13g2_inv_4 U5831 (.A(n172), .Y(N1110));
sg13g2_xnor2_1 U5832 (.A(keysched_new_key_o_131), .B(addroundkey_data_i_3), .Y(n40));
sg13g2_inv_4 U5833 (.A(n465), .Y(N817));
sg13g2_xnor2_1 U5834 (.A(key_i_104_), .B(addroundkey_data_i_40), .Y(n465));
sg13g2_inv_4 U5835 (.A(n209), .Y(N1073));
sg13g2_xnor2_1 U5836 (.A(keysched_new_key_o_168), .B(addroundkey_data_i_40), .Y(n77));
sg13g2_inv_4 U5837 (.A(n466), .Y(N816));
sg13g2_xnor2_1 U5838 (.A(key_i_105_), .B(addroundkey_data_i_41), .Y(n466));
sg13g2_inv_4 U5839 (.A(n210), .Y(N1072));
sg13g2_xnor2_1 U5840 (.A(keysched_new_key_o_169), .B(addroundkey_data_i_41), .Y(n78));
sg13g2_inv_4 U5841 (.A(n467), .Y(N815));
sg13g2_xnor2_1 U5842 (.A(key_i_106_), .B(addroundkey_data_i_42), .Y(n467));
sg13g2_inv_4 U5843 (.A(n211), .Y(N1071));
sg13g2_xnor2_1 U5844 (.A(keysched_new_key_o_170), .B(addroundkey_data_i_42), .Y(n79));
sg13g2_inv_4 U5845 (.A(n468), .Y(N814));
sg13g2_xnor2_1 U5846 (.A(key_i_107_), .B(addroundkey_data_i_43), .Y(n468));
sg13g2_inv_4 U5847 (.A(n212), .Y(N1070));
sg13g2_xnor2_1 U5848 (.A(keysched_new_key_o_171), .B(addroundkey_data_i_43), .Y(n80));
sg13g2_inv_4 U5849 (.A(n469), .Y(N813));
sg13g2_xnor2_1 U5850 (.A(key_i_108_), .B(addroundkey_data_i_44), .Y(n469));
sg13g2_inv_4 U5851 (.A(n213), .Y(N1069));
sg13g2_xnor2_1 U5852 (.A(keysched_new_key_o_172), .B(addroundkey_data_i_44), .Y(n81));
sg13g2_inv_4 U5853 (.A(n470), .Y(N812));
sg13g2_xnor2_1 U5854 (.A(key_i_109_), .B(addroundkey_data_i_45), .Y(n470));
sg13g2_inv_4 U5855 (.A(n214), .Y(N1068));
sg13g2_xnor2_1 U5856 (.A(keysched_new_key_o_173), .B(addroundkey_data_i_45), .Y(n82));
sg13g2_inv_4 U5857 (.A(n471), .Y(N811));
sg13g2_xnor2_1 U5858 (.A(key_i_110_), .B(addroundkey_data_i_46), .Y(n471));
sg13g2_inv_4 U5859 (.A(n215), .Y(N1067));
sg13g2_xnor2_1 U5860 (.A(keysched_new_key_o_174), .B(addroundkey_data_i_46), .Y(n83));
sg13g2_inv_4 U5861 (.A(n472), .Y(N810));
sg13g2_xnor2_1 U5862 (.A(key_i_111_), .B(addroundkey_data_i_47), .Y(n472));
sg13g2_inv_4 U5863 (.A(n216), .Y(N1066));
sg13g2_xnor2_1 U5864 (.A(keysched_new_key_o_175), .B(addroundkey_data_i_47), .Y(n84));
sg13g2_inv_4 U5865 (.A(n473), .Y(N809));
sg13g2_xnor2_1 U5866 (.A(key_i_112_), .B(addroundkey_data_i_48), .Y(n473));
sg13g2_inv_4 U5867 (.A(n217), .Y(N1065));
sg13g2_xnor2_1 U5868 (.A(keysched_new_key_o_176), .B(addroundkey_data_i_48), .Y(n85));
sg13g2_inv_4 U5869 (.A(n474), .Y(N808));
sg13g2_xnor2_1 U5870 (.A(key_i_113_), .B(addroundkey_data_i_49), .Y(n474));
sg13g2_inv_4 U5871 (.A(n218), .Y(N1064));
sg13g2_xnor2_1 U5872 (.A(keysched_new_key_o_177), .B(addroundkey_data_i_49), .Y(n86));
sg13g2_inv_4 U5873 (.A(n429), .Y(N853));
sg13g2_xnor2_1 U5874 (.A(key_i_68_), .B(addroundkey_data_i_4), .Y(n429));
sg13g2_inv_4 U5875 (.A(n173), .Y(N1109));
sg13g2_xnor2_1 U5876 (.A(keysched_new_key_o_132), .B(addroundkey_data_i_4), .Y(n41));
sg13g2_inv_4 U5877 (.A(n475), .Y(N807));
sg13g2_xnor2_1 U5878 (.A(key_i_114_), .B(addroundkey_data_i_50), .Y(n475));
sg13g2_inv_4 U5879 (.A(n219), .Y(N1063));
sg13g2_xnor2_1 U5880 (.A(keysched_new_key_o_178), .B(addroundkey_data_i_50), .Y(n87));
sg13g2_inv_4 U5881 (.A(n476), .Y(N806));
sg13g2_xnor2_1 U5882 (.A(key_i_115_), .B(addroundkey_data_i_51), .Y(n476));
sg13g2_inv_4 U5883 (.A(n220), .Y(N1062));
sg13g2_xnor2_1 U5884 (.A(keysched_new_key_o_179), .B(addroundkey_data_i_51), .Y(n88));
sg13g2_inv_4 U5885 (.A(n477), .Y(N805));
sg13g2_xnor2_1 U5886 (.A(key_i_116_), .B(addroundkey_data_i_52), .Y(n477));
sg13g2_inv_4 U5887 (.A(n221), .Y(N1061));
sg13g2_xnor2_1 U5888 (.A(keysched_new_key_o_180), .B(addroundkey_data_i_52), .Y(n89));
sg13g2_inv_4 U5889 (.A(n478), .Y(N804));
sg13g2_xnor2_1 U5890 (.A(key_i_117_), .B(addroundkey_data_i_53), .Y(n478));
sg13g2_inv_4 U5891 (.A(n222), .Y(N1060));
sg13g2_xnor2_1 U5892 (.A(keysched_new_key_o_181), .B(addroundkey_data_i_53), .Y(n90));
sg13g2_inv_4 U5893 (.A(n479), .Y(N803));
sg13g2_xnor2_1 U5894 (.A(key_i_118_), .B(addroundkey_data_i_54), .Y(n479));
sg13g2_inv_4 U5895 (.A(n223), .Y(N1059));
sg13g2_xnor2_1 U5896 (.A(keysched_new_key_o_182), .B(addroundkey_data_i_54), .Y(n91));
sg13g2_inv_4 U5897 (.A(n480), .Y(N802));
sg13g2_xnor2_1 U5898 (.A(key_i_119_), .B(addroundkey_data_i_55), .Y(n480));
sg13g2_inv_4 U5899 (.A(n224), .Y(N1058));
sg13g2_xnor2_1 U5900 (.A(keysched_new_key_o_183), .B(addroundkey_data_i_55), .Y(n92));
sg13g2_inv_4 U5901 (.A(n481), .Y(N801));
sg13g2_xnor2_1 U5902 (.A(key_i_120_), .B(addroundkey_data_i_56), .Y(n481));
sg13g2_inv_4 U5903 (.A(n225), .Y(N1057));
sg13g2_xnor2_1 U5904 (.A(keysched_new_key_o_184), .B(addroundkey_data_i_56), .Y(n93));
sg13g2_inv_4 U5905 (.A(n482), .Y(N800));
sg13g2_xnor2_1 U5906 (.A(key_i_121_), .B(addroundkey_data_i_57), .Y(n482));
sg13g2_inv_4 U5907 (.A(n226), .Y(N1056));
sg13g2_xnor2_1 U5908 (.A(keysched_new_key_o_185), .B(addroundkey_data_i_57), .Y(n94));
sg13g2_inv_4 U5909 (.A(n483), .Y(N799));
sg13g2_xnor2_1 U5910 (.A(key_i_122_), .B(addroundkey_data_i_58), .Y(n483));
sg13g2_inv_4 U5911 (.A(n227), .Y(N1055));
sg13g2_xnor2_1 U5912 (.A(keysched_new_key_o_186), .B(addroundkey_data_i_58), .Y(n95));
sg13g2_inv_4 U5913 (.A(n484), .Y(N798));
sg13g2_xnor2_1 U5914 (.A(key_i_123_), .B(addroundkey_data_i_59), .Y(n484));
sg13g2_inv_4 U5915 (.A(n228), .Y(N1054));
sg13g2_xnor2_1 U5916 (.A(keysched_new_key_o_187), .B(addroundkey_data_i_59), .Y(n96));
sg13g2_inv_4 U5917 (.A(n430), .Y(N852));
sg13g2_xnor2_1 U5918 (.A(key_i_69_), .B(addroundkey_data_i_5), .Y(n430));
sg13g2_inv_4 U5919 (.A(n174), .Y(N1108));
sg13g2_xnor2_1 U5920 (.A(keysched_new_key_o_133), .B(addroundkey_data_i_5), .Y(n42));
sg13g2_inv_4 U5921 (.A(n485), .Y(N797));
sg13g2_xnor2_1 U5922 (.A(key_i_124_), .B(addroundkey_data_i_60), .Y(n485));
sg13g2_inv_4 U5923 (.A(n229), .Y(N1053));
sg13g2_xnor2_1 U5924 (.A(keysched_new_key_o_188), .B(addroundkey_data_i_60), .Y(n97));
sg13g2_inv_4 U5925 (.A(n486), .Y(N796));
sg13g2_xnor2_1 U5926 (.A(key_i_125_), .B(addroundkey_data_i_61), .Y(n486));
sg13g2_inv_4 U5927 (.A(n230), .Y(N1052));
sg13g2_xnor2_1 U5928 (.A(keysched_new_key_o_189), .B(addroundkey_data_i_61), .Y(n98));
sg13g2_inv_4 U5929 (.A(n487), .Y(N795));
sg13g2_xnor2_1 U5930 (.A(key_i_126_), .B(addroundkey_data_i_62), .Y(n487));
sg13g2_inv_4 U5931 (.A(n231), .Y(N1051));
sg13g2_xnor2_1 U5932 (.A(keysched_new_key_o_190), .B(addroundkey_data_i_62), .Y(n99));
sg13g2_inv_4 U5933 (.A(n488), .Y(N794));
sg13g2_xnor2_1 U5934 (.A(key_i_127_), .B(addroundkey_data_i_63), .Y(n488));
sg13g2_inv_4 U5935 (.A(n232), .Y(N1050));
sg13g2_xnor2_1 U5936 (.A(keysched_new_key_o_191), .B(addroundkey_data_i_63), .Y(n100));
sg13g2_inv_4 U5937 (.A(n489), .Y(N793));
sg13g2_xnor2_1 U5938 (.A(key_i_128_), .B(addroundkey_data_i_64), .Y(n489));
sg13g2_inv_4 U5939 (.A(n233), .Y(N1049));
sg13g2_xnor2_1 U5940 (.A(N1342), .B(addroundkey_data_i_64), .Y(n101));
sg13g2_inv_4 U5941 (.A(n490), .Y(N792));
sg13g2_xnor2_1 U5942 (.A(key_i_129_), .B(addroundkey_data_i_65), .Y(n490));
sg13g2_inv_4 U5943 (.A(n234), .Y(N1048));
sg13g2_xnor2_1 U5944 (.A(N1343), .B(addroundkey_data_i_65), .Y(n102));
sg13g2_inv_4 U5945 (.A(n491), .Y(N791));
sg13g2_xnor2_1 U5946 (.A(key_i_130_), .B(addroundkey_data_i_66), .Y(n491));
sg13g2_inv_4 U5947 (.A(n235), .Y(N1047));
sg13g2_xnor2_1 U5948 (.A(N1344), .B(addroundkey_data_i_66), .Y(n103));
sg13g2_inv_4 U5949 (.A(n492), .Y(N790));
sg13g2_xnor2_1 U5950 (.A(key_i_131_), .B(addroundkey_data_i_67), .Y(n492));
sg13g2_inv_4 U5951 (.A(n236), .Y(N1046));
sg13g2_xnor2_1 U5952 (.A(N1345), .B(addroundkey_data_i_67), .Y(n104));
sg13g2_inv_4 U5953 (.A(n493), .Y(N789));
sg13g2_xnor2_1 U5954 (.A(key_i_132_), .B(addroundkey_data_i_68), .Y(n493));
sg13g2_inv_4 U5955 (.A(n237), .Y(N1045));
sg13g2_xnor2_1 U5956 (.A(N1346), .B(addroundkey_data_i_68), .Y(n105));
sg13g2_inv_4 U5957 (.A(n494), .Y(N788));
sg13g2_xnor2_1 U5958 (.A(key_i_133_), .B(addroundkey_data_i_69), .Y(n494));
sg13g2_inv_4 U5959 (.A(n238), .Y(N1044));
sg13g2_xnor2_1 U5960 (.A(N1347), .B(addroundkey_data_i_69), .Y(n106));
sg13g2_inv_4 U5961 (.A(n431), .Y(N851));
sg13g2_xnor2_1 U5962 (.A(key_i_70_), .B(addroundkey_data_i_6), .Y(n431));
sg13g2_inv_4 U5963 (.A(n175), .Y(N1107));
sg13g2_xnor2_1 U5964 (.A(keysched_new_key_o_134), .B(addroundkey_data_i_6), .Y(n43));
sg13g2_inv_4 U5965 (.A(n495), .Y(N787));
sg13g2_xnor2_1 U5966 (.A(key_i_134_), .B(addroundkey_data_i_70), .Y(n495));
sg13g2_inv_4 U5967 (.A(n239), .Y(N1043));
sg13g2_xnor2_1 U5968 (.A(N1348), .B(addroundkey_data_i_70), .Y(n107));
sg13g2_inv_4 U5969 (.A(n496), .Y(N786));
sg13g2_xnor2_1 U5970 (.A(key_i_135_), .B(addroundkey_data_i_71), .Y(n496));
sg13g2_inv_4 U5971 (.A(n240), .Y(N1042));
sg13g2_xnor2_1 U5972 (.A(N1349), .B(addroundkey_data_i_71), .Y(n108));
sg13g2_inv_4 U5973 (.A(n497), .Y(N785));
sg13g2_xnor2_1 U5974 (.A(key_i_136_), .B(addroundkey_data_i_72), .Y(n497));
sg13g2_inv_4 U5975 (.A(n241), .Y(N1041));
sg13g2_xnor2_1 U5976 (.A(N1350), .B(addroundkey_data_i_72), .Y(n109));
sg13g2_inv_4 U5977 (.A(n499), .Y(N783));
sg13g2_xnor2_1 U5978 (.A(key_i_138_), .B(addroundkey_data_i_74), .Y(n499));
sg13g2_inv_4 U5979 (.A(n243), .Y(N1039));
sg13g2_xnor2_1 U5980 (.A(N1352), .B(addroundkey_data_i_74), .Y(n111));
sg13g2_inv_4 U5981 (.A(n500), .Y(N782));
sg13g2_xnor2_1 U5982 (.A(key_i_139_), .B(addroundkey_data_i_75), .Y(n500));
sg13g2_inv_4 U5983 (.A(n244), .Y(N1038));
sg13g2_xnor2_1 U5984 (.A(N1353), .B(addroundkey_data_i_75), .Y(n112));
sg13g2_inv_4 U5985 (.A(n501), .Y(N781));
sg13g2_xnor2_1 U5986 (.A(key_i_140_), .B(addroundkey_data_i_76), .Y(n501));
sg13g2_inv_4 U5987 (.A(n245), .Y(N1037));
sg13g2_xnor2_1 U5988 (.A(N1354), .B(addroundkey_data_i_76), .Y(n113));
sg13g2_inv_4 U5989 (.A(n502), .Y(N780));
sg13g2_xnor2_1 U5990 (.A(key_i_141_), .B(addroundkey_data_i_77), .Y(n502));
sg13g2_inv_4 U5991 (.A(n246), .Y(N1036));
sg13g2_xnor2_1 U5992 (.A(N1355), .B(addroundkey_data_i_77), .Y(n114));
sg13g2_inv_4 U5993 (.A(n503), .Y(N779));
sg13g2_xnor2_1 U5994 (.A(key_i_142_), .B(addroundkey_data_i_78), .Y(n503));
sg13g2_inv_4 U5995 (.A(n247), .Y(N1035));
sg13g2_xnor2_1 U5996 (.A(N1356), .B(addroundkey_data_i_78), .Y(n115));
sg13g2_inv_4 U5997 (.A(n504), .Y(N778));
sg13g2_xnor2_1 U5998 (.A(key_i_143_), .B(addroundkey_data_i_79), .Y(n504));
sg13g2_inv_4 U5999 (.A(n248), .Y(N1034));
sg13g2_xnor2_1 U6000 (.A(N1357), .B(addroundkey_data_i_79), .Y(n116));
sg13g2_inv_4 U6001 (.A(n432), .Y(N850));
sg13g2_xnor2_1 U6002 (.A(key_i_71_), .B(addroundkey_data_i_7), .Y(n432));
sg13g2_inv_4 U6003 (.A(n176), .Y(N1106));
sg13g2_xnor2_1 U6004 (.A(keysched_new_key_o_135), .B(addroundkey_data_i_7), .Y(n44));
sg13g2_inv_4 U6005 (.A(n505), .Y(N777));
sg13g2_xnor2_1 U6006 (.A(key_i_144_), .B(addroundkey_data_i_80), .Y(n505));
sg13g2_inv_4 U6007 (.A(n249), .Y(N1033));
sg13g2_xnor2_1 U6008 (.A(N1358), .B(addroundkey_data_i_80), .Y(n117));
sg13g2_inv_4 U6009 (.A(n506), .Y(N776));
sg13g2_xnor2_1 U6010 (.A(key_i_145_), .B(addroundkey_data_i_81), .Y(n506));
sg13g2_inv_4 U6011 (.A(n250), .Y(N1032));
sg13g2_xnor2_1 U6012 (.A(N1359), .B(addroundkey_data_i_81), .Y(n118));
sg13g2_inv_4 U6013 (.A(n507), .Y(N775));
sg13g2_xnor2_1 U6014 (.A(key_i_146_), .B(addroundkey_data_i_82), .Y(n507));
sg13g2_inv_4 U6015 (.A(n251), .Y(N1031));
sg13g2_xnor2_1 U6016 (.A(N1360), .B(addroundkey_data_i_82), .Y(n119));
sg13g2_inv_4 U6017 (.A(n508), .Y(N774));
sg13g2_xnor2_1 U6018 (.A(key_i_147_), .B(addroundkey_data_i_83), .Y(n508));
sg13g2_inv_4 U6019 (.A(n252), .Y(N1030));
sg13g2_xnor2_1 U6020 (.A(N1361), .B(addroundkey_data_i_83), .Y(n120));
sg13g2_inv_4 U6021 (.A(n509), .Y(N773));
sg13g2_xnor2_1 U6022 (.A(key_i_148_), .B(addroundkey_data_i_84), .Y(n509));
sg13g2_inv_4 U6023 (.A(n253), .Y(N1029));
sg13g2_xnor2_1 U6024 (.A(N1362), .B(addroundkey_data_i_84), .Y(n121));
sg13g2_inv_4 U6025 (.A(n510), .Y(N772));
sg13g2_xnor2_1 U6026 (.A(key_i_149_), .B(addroundkey_data_i_85), .Y(n510));
sg13g2_inv_4 U6027 (.A(n254), .Y(N1028));
sg13g2_xnor2_1 U6028 (.A(N1363), .B(addroundkey_data_i_85), .Y(n122));
sg13g2_inv_4 U6029 (.A(n511), .Y(N771));
sg13g2_xnor2_1 U6030 (.A(key_i_150_), .B(addroundkey_data_i_86), .Y(n511));
sg13g2_inv_4 U6031 (.A(n255), .Y(N1027));
sg13g2_xnor2_1 U6032 (.A(N1364), .B(addroundkey_data_i_86), .Y(n123));
sg13g2_inv_4 U6033 (.A(n512), .Y(N770));
sg13g2_xnor2_1 U6034 (.A(key_i_151_), .B(addroundkey_data_i_87), .Y(n512));
sg13g2_inv_4 U6035 (.A(n256), .Y(N1026));
sg13g2_xnor2_1 U6036 (.A(N1365), .B(addroundkey_data_i_87), .Y(n124));
sg13g2_inv_4 U6037 (.A(n513), .Y(N769));
sg13g2_xnor2_1 U6038 (.A(key_i_152_), .B(addroundkey_data_i_88), .Y(n513));
sg13g2_inv_4 U6039 (.A(n257), .Y(N1025));
sg13g2_xnor2_1 U6040 (.A(N1366), .B(addroundkey_data_i_88), .Y(n125));
sg13g2_inv_4 U6041 (.A(n514), .Y(N768));
sg13g2_xnor2_1 U6042 (.A(key_i_153_), .B(addroundkey_data_i_89), .Y(n514));
sg13g2_inv_4 U6043 (.A(n258), .Y(N1024));
sg13g2_xnor2_1 U6044 (.A(N1367), .B(addroundkey_data_i_89), .Y(n126));
sg13g2_inv_4 U6045 (.A(n433), .Y(N849));
sg13g2_xnor2_1 U6046 (.A(key_i_72_), .B(addroundkey_data_i_8), .Y(n433));
sg13g2_inv_4 U6047 (.A(n177), .Y(N1105));
sg13g2_xnor2_1 U6048 (.A(keysched_new_key_o_136), .B(addroundkey_data_i_8), .Y(n45));
sg13g2_inv_4 U6049 (.A(n515), .Y(N767));
sg13g2_xnor2_1 U6050 (.A(key_i_154_), .B(addroundkey_data_i_90), .Y(n515));
sg13g2_inv_4 U6051 (.A(n259), .Y(N1023));
sg13g2_xnor2_1 U6052 (.A(N1368), .B(addroundkey_data_i_90), .Y(n127));
sg13g2_inv_4 U6053 (.A(n516), .Y(N766));
sg13g2_xnor2_1 U6054 (.A(key_i_155_), .B(addroundkey_data_i_91), .Y(n516));
sg13g2_inv_4 U6055 (.A(n260), .Y(N1022));
sg13g2_xnor2_1 U6056 (.A(N1369), .B(addroundkey_data_i_91), .Y(n128));
sg13g2_inv_4 U6057 (.A(n517), .Y(N765));
sg13g2_xnor2_1 U6058 (.A(key_i_156_), .B(addroundkey_data_i_92), .Y(n517));
sg13g2_inv_4 U6059 (.A(n261), .Y(N1021));
sg13g2_xnor2_1 U6060 (.A(N1370), .B(addroundkey_data_i_92), .Y(n129));
sg13g2_inv_4 U6061 (.A(n518), .Y(N764));
sg13g2_xnor2_1 U6062 (.A(key_i_157_), .B(addroundkey_data_i_93), .Y(n518));
sg13g2_inv_4 U6063 (.A(n262), .Y(N1020));
sg13g2_xnor2_1 U6064 (.A(N1371), .B(addroundkey_data_i_93), .Y(n130));
sg13g2_inv_4 U6065 (.A(n519), .Y(N763));
sg13g2_xnor2_1 U6066 (.A(key_i_158_), .B(addroundkey_data_i_94), .Y(n519));
sg13g2_inv_4 U6067 (.A(n263), .Y(N1019));
sg13g2_xnor2_1 U6068 (.A(N1372), .B(addroundkey_data_i_94), .Y(n131));
sg13g2_inv_4 U6069 (.A(n520), .Y(N762));
sg13g2_xnor2_1 U6070 (.A(key_i_159_), .B(addroundkey_data_i_95), .Y(n520));
sg13g2_inv_4 U6071 (.A(n264), .Y(N1018));
sg13g2_xnor2_1 U6072 (.A(N1373), .B(addroundkey_data_i_95), .Y(n132));
sg13g2_inv_4 U6073 (.A(n521), .Y(N761));
sg13g2_xnor2_1 U6074 (.A(key_i_160_), .B(addroundkey_data_i_96), .Y(n521));
sg13g2_inv_4 U6075 (.A(n265), .Y(N1017));
sg13g2_xnor2_1 U6076 (.A(N1374), .B(addroundkey_data_i_96), .Y(n133));
sg13g2_inv_4 U6077 (.A(n522), .Y(N760));
sg13g2_xnor2_1 U6078 (.A(key_i_161_), .B(addroundkey_data_i_97), .Y(n522));
sg13g2_inv_4 U6079 (.A(n266), .Y(N1016));
sg13g2_xnor2_1 U6080 (.A(N1375), .B(addroundkey_data_i_97), .Y(n134));
sg13g2_inv_4 U6081 (.A(n523), .Y(N759));
sg13g2_xnor2_1 U6082 (.A(key_i_162_), .B(addroundkey_data_i_98), .Y(n523));
sg13g2_inv_4 U6083 (.A(n267), .Y(N1015));
sg13g2_xnor2_1 U6084 (.A(N1376), .B(addroundkey_data_i_98), .Y(n135));
sg13g2_inv_4 U6085 (.A(n524), .Y(N758));
sg13g2_xnor2_1 U6086 (.A(key_i_163_), .B(addroundkey_data_i_99), .Y(n524));
sg13g2_inv_4 U6087 (.A(n268), .Y(N1014));
sg13g2_xnor2_1 U6088 (.A(N1377), .B(addroundkey_data_i_99), .Y(n136));
sg13g2_inv_4 U6089 (.A(n434), .Y(N848));
sg13g2_xnor2_1 U6090 (.A(key_i_73_), .B(addroundkey_data_i_9), .Y(n434));
sg13g2_inv_4 U6091 (.A(n178), .Y(N1104));
sg13g2_xnor2_1 U6092 (.A(keysched_new_key_o_137), .B(addroundkey_data_i_9), .Y(n46));
sg13g2_inv_4 U6093 (.A(n425), .Y(N857));
sg13g2_xnor2_1 U6094 (.A(key_i_64_), .B(addroundkey_data_i_0), .Y(n425));
sg13g2_inv_4 U6095 (.A(n169), .Y(N1113));
sg13g2_xnor2_1 U6096 (.A(keysched_new_key_o_128), .B(addroundkey_data_i_0), .Y(n37));
sg13g2_inv_4 U6097 (.A(n498), .Y(N784));
sg13g2_xnor2_1 U6098 (.A(key_i_137_), .B(addroundkey_data_i_73), .Y(n498));
sg13g2_inv_4 U6099 (.A(n242), .Y(N1040));
sg13g2_xnor2_1 U6100 (.A(N1351), .B(addroundkey_data_i_73), .Y(n110));
sg13g2_inv_4 U6101 (.A(n3701), .Y(N1119));
sg13g2_inv_4 U6102 (.A(decrypt_i), .Y(N29));
sg13g2_xnor2_1 U6108 (.A(keysched_new_key_o_164), .B(addroundkey_data_i_100), .Y(n397));
sg13g2_xnor2_1 U6110 (.A(keysched_new_key_o_165), .B(addroundkey_data_i_101), .Y(n398));
sg13g2_xnor2_1 U6112 (.A(keysched_new_key_o_166), .B(addroundkey_data_i_102), .Y(n399));
sg13g2_xnor2_1 U6114 (.A(keysched_new_key_o_167), .B(addroundkey_data_i_103), .Y(n400));
sg13g2_xnor2_1 U6116 (.A(keysched_new_key_o_168), .B(addroundkey_data_i_104), .Y(n401));
sg13g2_xnor2_1 U6118 (.A(keysched_new_key_o_169), .B(addroundkey_data_i_105), .Y(n402));
sg13g2_xnor2_1 U6120 (.A(keysched_new_key_o_170), .B(addroundkey_data_i_106), .Y(n403));
sg13g2_xnor2_1 U6122 (.A(keysched_new_key_o_171), .B(addroundkey_data_i_107), .Y(n404));
sg13g2_xnor2_1 U6124 (.A(keysched_new_key_o_172), .B(addroundkey_data_i_108), .Y(n405));
sg13g2_xnor2_1 U6126 (.A(keysched_new_key_o_173), .B(addroundkey_data_i_109), .Y(n406));
sg13g2_xnor2_1 U6128 (.A(keysched_new_key_o_74), .B(addroundkey_data_i_10), .Y(n307));
sg13g2_xnor2_1 U6130 (.A(keysched_new_key_o_174), .B(addroundkey_data_i_110), .Y(n407));
sg13g2_xnor2_1 U6132 (.A(keysched_new_key_o_175), .B(addroundkey_data_i_111), .Y(n408));
sg13g2_xnor2_1 U6134 (.A(keysched_new_key_o_176), .B(addroundkey_data_i_112), .Y(n409));
sg13g2_xnor2_1 U6136 (.A(keysched_new_key_o_177), .B(addroundkey_data_i_113), .Y(n410));
sg13g2_xnor2_1 U6138 (.A(keysched_new_key_o_178), .B(addroundkey_data_i_114), .Y(n411));
sg13g2_xnor2_1 U6140 (.A(keysched_new_key_o_179), .B(addroundkey_data_i_115), .Y(n412));
sg13g2_xnor2_1 U6142 (.A(keysched_new_key_o_180), .B(addroundkey_data_i_116), .Y(n413));
sg13g2_xnor2_1 U6144 (.A(keysched_new_key_o_181), .B(addroundkey_data_i_117), .Y(n414));
sg13g2_xnor2_1 U6146 (.A(keysched_new_key_o_182), .B(addroundkey_data_i_118), .Y(n415));
sg13g2_xnor2_1 U6148 (.A(keysched_new_key_o_183), .B(addroundkey_data_i_119), .Y(n416));
sg13g2_xnor2_1 U6150 (.A(keysched_new_key_o_75), .B(addroundkey_data_i_11), .Y(n308));
sg13g2_xnor2_1 U6152 (.A(keysched_new_key_o_184), .B(addroundkey_data_i_120), .Y(n417));
sg13g2_xnor2_1 U6154 (.A(keysched_new_key_o_185), .B(addroundkey_data_i_121), .Y(n418));
sg13g2_xnor2_1 U6156 (.A(keysched_new_key_o_186), .B(addroundkey_data_i_122), .Y(n419));
sg13g2_xnor2_1 U6158 (.A(keysched_new_key_o_187), .B(addroundkey_data_i_123), .Y(n420));
sg13g2_xnor2_1 U6160 (.A(keysched_new_key_o_188), .B(addroundkey_data_i_124), .Y(n421));
sg13g2_xnor2_1 U6162 (.A(keysched_new_key_o_189), .B(addroundkey_data_i_125), .Y(n422));
sg13g2_xnor2_1 U6164 (.A(keysched_new_key_o_190), .B(addroundkey_data_i_126), .Y(n423));
sg13g2_xnor2_1 U6166 (.A(keysched_new_key_o_191), .B(addroundkey_data_i_127), .Y(n424));
sg13g2_xnor2_1 U6168 (.A(keysched_new_key_o_76), .B(addroundkey_data_i_12), .Y(n309));
sg13g2_xnor2_1 U6170 (.A(keysched_new_key_o_77), .B(addroundkey_data_i_13), .Y(n310));
sg13g2_xnor2_1 U6172 (.A(keysched_new_key_o_78), .B(addroundkey_data_i_14), .Y(n311));
sg13g2_xnor2_1 U6174 (.A(keysched_new_key_o_79), .B(addroundkey_data_i_15), .Y(n312));
sg13g2_xnor2_1 U6176 (.A(keysched_new_key_o_80), .B(addroundkey_data_i_16), .Y(n313));
sg13g2_xnor2_1 U6178 (.A(keysched_new_key_o_81), .B(addroundkey_data_i_17), .Y(n314));
sg13g2_xnor2_1 U6180 (.A(keysched_new_key_o_82), .B(addroundkey_data_i_18), .Y(n315));
sg13g2_xnor2_1 U6182 (.A(keysched_new_key_o_83), .B(addroundkey_data_i_19), .Y(n316));
sg13g2_xnor2_1 U6184 (.A(keysched_new_key_o_65), .B(addroundkey_data_i_1), .Y(n298));
sg13g2_xnor2_1 U6186 (.A(keysched_new_key_o_84), .B(addroundkey_data_i_20), .Y(n317));
sg13g2_xnor2_1 U6188 (.A(keysched_new_key_o_85), .B(addroundkey_data_i_21), .Y(n318));
sg13g2_xnor2_1 U6190 (.A(keysched_new_key_o_86), .B(addroundkey_data_i_22), .Y(n319));
sg13g2_xnor2_1 U6192 (.A(keysched_new_key_o_87), .B(addroundkey_data_i_23), .Y(n320));
sg13g2_xnor2_1 U6194 (.A(keysched_new_key_o_88), .B(addroundkey_data_i_24), .Y(n321));
sg13g2_xnor2_1 U6196 (.A(keysched_new_key_o_89), .B(addroundkey_data_i_25), .Y(n322));
sg13g2_xnor2_1 U6198 (.A(keysched_new_key_o_90), .B(addroundkey_data_i_26), .Y(n323));
sg13g2_xnor2_1 U6200 (.A(keysched_new_key_o_91), .B(addroundkey_data_i_27), .Y(n324));
sg13g2_xnor2_1 U6202 (.A(keysched_new_key_o_92), .B(addroundkey_data_i_28), .Y(n325));
sg13g2_xnor2_1 U6204 (.A(keysched_new_key_o_93), .B(addroundkey_data_i_29), .Y(n326));
sg13g2_xnor2_1 U6206 (.A(keysched_new_key_o_66), .B(addroundkey_data_i_2), .Y(n299));
sg13g2_xnor2_1 U6208 (.A(keysched_new_key_o_94), .B(addroundkey_data_i_30), .Y(n327));
sg13g2_xnor2_1 U6210 (.A(keysched_new_key_o_95), .B(addroundkey_data_i_31), .Y(n328));
sg13g2_xnor2_1 U6212 (.A(keysched_new_key_o_96), .B(addroundkey_data_i_32), .Y(n329));
sg13g2_xnor2_1 U6214 (.A(keysched_new_key_o_97), .B(addroundkey_data_i_33), .Y(n330));
sg13g2_xnor2_1 U6216 (.A(keysched_new_key_o_98), .B(addroundkey_data_i_34), .Y(n331));
sg13g2_xnor2_1 U6218 (.A(keysched_new_key_o_99), .B(addroundkey_data_i_35), .Y(n332));
sg13g2_xnor2_1 U6220 (.A(keysched_new_key_o_100), .B(addroundkey_data_i_36), .Y(n333));
sg13g2_xnor2_1 U6222 (.A(keysched_new_key_o_101), .B(addroundkey_data_i_37), .Y(n334));
sg13g2_xnor2_1 U6224 (.A(keysched_new_key_o_102), .B(addroundkey_data_i_38), .Y(n335));
sg13g2_xnor2_1 U6226 (.A(keysched_new_key_o_103), .B(addroundkey_data_i_39), .Y(n336));
sg13g2_xnor2_1 U6228 (.A(keysched_new_key_o_67), .B(addroundkey_data_i_3), .Y(n300));
sg13g2_xnor2_1 U6230 (.A(keysched_new_key_o_104), .B(addroundkey_data_i_40), .Y(n337));
sg13g2_xnor2_1 U6232 (.A(keysched_new_key_o_105), .B(addroundkey_data_i_41), .Y(n338));
sg13g2_xnor2_1 U6234 (.A(keysched_new_key_o_106), .B(addroundkey_data_i_42), .Y(n339));
sg13g2_xnor2_1 U6236 (.A(keysched_new_key_o_107), .B(addroundkey_data_i_43), .Y(n340));
sg13g2_xnor2_1 U6238 (.A(keysched_new_key_o_108), .B(addroundkey_data_i_44), .Y(n341));
sg13g2_xnor2_1 U6240 (.A(keysched_new_key_o_109), .B(addroundkey_data_i_45), .Y(n342));
sg13g2_xnor2_1 U6242 (.A(keysched_new_key_o_110), .B(addroundkey_data_i_46), .Y(n343));
sg13g2_xnor2_1 U6244 (.A(keysched_new_key_o_111), .B(addroundkey_data_i_47), .Y(n344));
sg13g2_xnor2_1 U6246 (.A(keysched_new_key_o_112), .B(addroundkey_data_i_48), .Y(n345));
sg13g2_xnor2_1 U6248 (.A(keysched_new_key_o_113), .B(addroundkey_data_i_49), .Y(n346));
sg13g2_xnor2_1 U6250 (.A(keysched_new_key_o_68), .B(addroundkey_data_i_4), .Y(n301));
sg13g2_xnor2_1 U6252 (.A(keysched_new_key_o_114), .B(addroundkey_data_i_50), .Y(n347));
sg13g2_xnor2_1 U6254 (.A(keysched_new_key_o_115), .B(addroundkey_data_i_51), .Y(n348));
sg13g2_xnor2_1 U6256 (.A(keysched_new_key_o_116), .B(addroundkey_data_i_52), .Y(n349));
sg13g2_xnor2_1 U6258 (.A(keysched_new_key_o_117), .B(addroundkey_data_i_53), .Y(n350));
sg13g2_xnor2_1 U6260 (.A(keysched_new_key_o_118), .B(addroundkey_data_i_54), .Y(n351));
sg13g2_xnor2_1 U6262 (.A(keysched_new_key_o_119), .B(addroundkey_data_i_55), .Y(n352));
sg13g2_xnor2_1 U6264 (.A(keysched_new_key_o_120), .B(addroundkey_data_i_56), .Y(n353));
sg13g2_xnor2_1 U6266 (.A(keysched_new_key_o_121), .B(addroundkey_data_i_57), .Y(n354));
sg13g2_xnor2_1 U6268 (.A(keysched_new_key_o_122), .B(addroundkey_data_i_58), .Y(n355));
sg13g2_xnor2_1 U6270 (.A(keysched_new_key_o_123), .B(addroundkey_data_i_59), .Y(n356));
sg13g2_xnor2_1 U6272 (.A(keysched_new_key_o_69), .B(addroundkey_data_i_5), .Y(n302));
sg13g2_xnor2_1 U6274 (.A(keysched_new_key_o_124), .B(addroundkey_data_i_60), .Y(n357));
sg13g2_xnor2_1 U6276 (.A(keysched_new_key_o_125), .B(addroundkey_data_i_61), .Y(n358));
sg13g2_xnor2_1 U6278 (.A(keysched_new_key_o_126), .B(addroundkey_data_i_62), .Y(n359));
sg13g2_xnor2_1 U6280 (.A(keysched_new_key_o_127), .B(addroundkey_data_i_63), .Y(n360));
sg13g2_xnor2_1 U6282 (.A(keysched_new_key_o_128), .B(addroundkey_data_i_64), .Y(n361));
sg13g2_xnor2_1 U6284 (.A(keysched_new_key_o_129), .B(addroundkey_data_i_65), .Y(n362));
sg13g2_xnor2_1 U6286 (.A(keysched_new_key_o_130), .B(addroundkey_data_i_66), .Y(n363));
sg13g2_xnor2_1 U6288 (.A(keysched_new_key_o_131), .B(addroundkey_data_i_67), .Y(n364));
sg13g2_xnor2_1 U6290 (.A(keysched_new_key_o_132), .B(addroundkey_data_i_68), .Y(n365));
sg13g2_xnor2_1 U6292 (.A(keysched_new_key_o_133), .B(addroundkey_data_i_69), .Y(n366));
sg13g2_xnor2_1 U6294 (.A(keysched_new_key_o_70), .B(addroundkey_data_i_6), .Y(n303));
sg13g2_xnor2_1 U6296 (.A(keysched_new_key_o_134), .B(addroundkey_data_i_70), .Y(n367));
sg13g2_xnor2_1 U6298 (.A(keysched_new_key_o_135), .B(addroundkey_data_i_71), .Y(n368));
sg13g2_xnor2_1 U6300 (.A(keysched_new_key_o_136), .B(addroundkey_data_i_72), .Y(n369));
sg13g2_xnor2_1 U6302 (.A(keysched_new_key_o_138), .B(addroundkey_data_i_74), .Y(n371));
sg13g2_xnor2_1 U6304 (.A(keysched_new_key_o_139), .B(addroundkey_data_i_75), .Y(n372));
sg13g2_xnor2_1 U6306 (.A(keysched_new_key_o_140), .B(addroundkey_data_i_76), .Y(n373));
sg13g2_xnor2_1 U6308 (.A(keysched_new_key_o_141), .B(addroundkey_data_i_77), .Y(n374));
sg13g2_xnor2_1 U6310 (.A(keysched_new_key_o_142), .B(addroundkey_data_i_78), .Y(n375));
sg13g2_xnor2_1 U6312 (.A(keysched_new_key_o_143), .B(addroundkey_data_i_79), .Y(n376));
sg13g2_xnor2_1 U6314 (.A(keysched_new_key_o_71), .B(addroundkey_data_i_7), .Y(n304));
sg13g2_xnor2_1 U6316 (.A(keysched_new_key_o_144), .B(addroundkey_data_i_80), .Y(n377));
sg13g2_xnor2_1 U6318 (.A(keysched_new_key_o_145), .B(addroundkey_data_i_81), .Y(n378));
sg13g2_xnor2_1 U6320 (.A(keysched_new_key_o_146), .B(addroundkey_data_i_82), .Y(n379));
sg13g2_xnor2_1 U6322 (.A(keysched_new_key_o_147), .B(addroundkey_data_i_83), .Y(n380));
sg13g2_xnor2_1 U6324 (.A(keysched_new_key_o_148), .B(addroundkey_data_i_84), .Y(n381));
sg13g2_xnor2_1 U6326 (.A(keysched_new_key_o_149), .B(addroundkey_data_i_85), .Y(n382));
sg13g2_xnor2_1 U6328 (.A(keysched_new_key_o_150), .B(addroundkey_data_i_86), .Y(n383));
sg13g2_xnor2_1 U6330 (.A(keysched_new_key_o_151), .B(addroundkey_data_i_87), .Y(n384));
sg13g2_xnor2_1 U6332 (.A(keysched_new_key_o_152), .B(addroundkey_data_i_88), .Y(n385));
sg13g2_xnor2_1 U6334 (.A(keysched_new_key_o_153), .B(addroundkey_data_i_89), .Y(n386));
sg13g2_xnor2_1 U6336 (.A(keysched_new_key_o_72), .B(addroundkey_data_i_8), .Y(n305));
sg13g2_xnor2_1 U6338 (.A(keysched_new_key_o_154), .B(addroundkey_data_i_90), .Y(n387));
sg13g2_xnor2_1 U6340 (.A(keysched_new_key_o_155), .B(addroundkey_data_i_91), .Y(n388));
sg13g2_xnor2_1 U6342 (.A(keysched_new_key_o_156), .B(addroundkey_data_i_92), .Y(n389));
sg13g2_xnor2_1 U6344 (.A(keysched_new_key_o_157), .B(addroundkey_data_i_93), .Y(n390));
sg13g2_xnor2_1 U6346 (.A(keysched_new_key_o_158), .B(addroundkey_data_i_94), .Y(n391));
sg13g2_xnor2_1 U6348 (.A(keysched_new_key_o_159), .B(addroundkey_data_i_95), .Y(n392));
sg13g2_xnor2_1 U6350 (.A(keysched_new_key_o_160), .B(addroundkey_data_i_96), .Y(n393));
sg13g2_xnor2_1 U6352 (.A(keysched_new_key_o_161), .B(addroundkey_data_i_97), .Y(n394));
sg13g2_xnor2_1 U6354 (.A(keysched_new_key_o_162), .B(addroundkey_data_i_98), .Y(n395));
sg13g2_xnor2_1 U6356 (.A(keysched_new_key_o_163), .B(addroundkey_data_i_99), .Y(n396));
sg13g2_xnor2_1 U6358 (.A(keysched_new_key_o_73), .B(addroundkey_data_i_9), .Y(n306));
sg13g2_xnor2_1 U6426 (.A(keysched_new_key_o_64), .B(addroundkey_data_i_0), .Y(n297));
sg13g2_xnor2_1 U6427 (.A(keysched_new_key_o_137), .B(addroundkey_data_i_73), .Y(n370));
sg13g2_buf_8 U6429 (.A(n4266), .X(n4325));
sg13g2_buf_8 U6430 (.A(n4266), .X(n4326));
sg13g2_buf_8 U6431 (.A(n4266), .X(n4327));
sg13g2_buf_8 U6432 (.A(n4162), .X(n4328));
sg13g2_buf_8 U6433 (.A(n4266), .X(n4329));
sg13g2_buf_8 U6434 (.A(n4162), .X(n4330));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_0_ (.CLK(clk), .D(n4128), .Q(data_o_0_), .Q_N(n1773), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_1_ (.CLK(clk), .D(n4127), .Q(data_o_1_), .Q_N(n1578), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_2_ (.CLK(clk), .D(n4126), .Q(data_o_2_), .Q_N(n1523), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_3_ (.CLK(clk), .D(n4125), .Q(data_o_3_), .Q_N(n1468), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_4_ (.CLK(clk), .D(n4124), .Q(data_o_4_), .Q_N(n1413), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_5_ (.CLK(clk), .D(n4123), .Q(data_o_5_), .Q_N(n1358), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_6_ (.CLK(clk), .D(n4122), .Q(data_o_6_), .Q_N(n1303), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_7_ (.CLK(clk), .D(n4121), .Q(data_o_7_), .Q_N(n1248), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_8_ (.CLK(clk), .D(n4120), .Q(data_o_8_), .Q_N(n1193), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_9_ (.CLK(clk), .D(n4119), .Q(data_o_9_), .Q_N(n1136), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_10_ (.CLK(clk), .D(n4118), .Q(data_o_10_), .Q_N(n1718), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_11_ (.CLK(clk), .D(n4117), .Q(data_o_11_), .Q_N(n1663), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_12_ (.CLK(clk), .D(n4116), .Q(data_o_12_), .Q_N(n1618), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_13_ (.CLK(clk), .D(n4115), .Q(data_o_13_), .Q_N(n1613), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_14_ (.CLK(clk), .D(n4114), .Q(data_o_14_), .Q_N(n1608), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_15_ (.CLK(clk), .D(n4113), .Q(data_o_15_), .Q_N(n1603), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_16_ (.CLK(clk), .D(n4112), .Q(data_o_16_), .Q_N(n1598), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_17_ (.CLK(clk), .D(n4111), .Q(data_o_17_), .Q_N(n1593), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_18_ (.CLK(clk), .D(n4110), .Q(data_o_18_), .Q_N(n1588), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_19_ (.CLK(clk), .D(n4109), .Q(data_o_19_), .Q_N(n1583), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_20_ (.CLK(clk), .D(n4108), .Q(data_o_20_), .Q_N(n1573), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_21_ (.CLK(clk), .D(n4107), .Q(data_o_21_), .Q_N(n1568), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_22_ (.CLK(clk), .D(n4106), .Q(data_o_22_), .Q_N(n1563), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_23_ (.CLK(clk), .D(n4105), .Q(data_o_23_), .Q_N(n1558), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_24_ (.CLK(clk), .D(n4104), .Q(data_o_24_), .Q_N(n1553), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_25_ (.CLK(clk), .D(n4103), .Q(data_o_25_), .Q_N(n1548), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_26_ (.CLK(clk), .D(n4102), .Q(data_o_26_), .Q_N(n1543), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_27_ (.CLK(clk), .D(n4101), .Q(data_o_27_), .Q_N(n1538), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_28_ (.CLK(clk), .D(n4100), .Q(data_o_28_), .Q_N(n1533), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_29_ (.CLK(clk), .D(n4099), .Q(data_o_29_), .Q_N(n1528), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_30_ (.CLK(clk), .D(n4098), .Q(data_o_30_), .Q_N(n1518), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_31_ (.CLK(clk), .D(n4097), .Q(data_o_31_), .Q_N(n1513), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_32_ (.CLK(clk), .D(n4096), .Q(data_o_32_), .Q_N(n1508), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_33_ (.CLK(clk), .D(n4095), .Q(data_o_33_), .Q_N(n1503), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_34_ (.CLK(clk), .D(n4094), .Q(data_o_34_), .Q_N(n1498), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_35_ (.CLK(clk), .D(n4093), .Q(data_o_35_), .Q_N(n1493), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_36_ (.CLK(clk), .D(n4092), .Q(data_o_36_), .Q_N(n1488), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_37_ (.CLK(clk), .D(n4091), .Q(data_o_37_), .Q_N(n1483), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_38_ (.CLK(clk), .D(n4090), .Q(data_o_38_), .Q_N(n1478), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_39_ (.CLK(clk), .D(n4089), .Q(data_o_39_), .Q_N(n1473), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_40_ (.CLK(clk), .D(n4088), .Q(data_o_40_), .Q_N(n1463), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_41_ (.CLK(clk), .D(n4087), .Q(data_o_41_), .Q_N(n1458), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_42_ (.CLK(clk), .D(n4086), .Q(data_o_42_), .Q_N(n1453), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_43_ (.CLK(clk), .D(n4085), .Q(data_o_43_), .Q_N(n1448), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_44_ (.CLK(clk), .D(n4084), .Q(data_o_44_), .Q_N(n1443), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_45_ (.CLK(clk), .D(n4083), .Q(data_o_45_), .Q_N(n1438), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_46_ (.CLK(clk), .D(n4082), .Q(data_o_46_), .Q_N(n1433), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_47_ (.CLK(clk), .D(n4081), .Q(data_o_47_), .Q_N(n1428), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_48_ (.CLK(clk), .D(n4080), .Q(data_o_48_), .Q_N(n1423), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_49_ (.CLK(clk), .D(n4079), .Q(data_o_49_), .Q_N(n1418), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_50_ (.CLK(clk), .D(n4078), .Q(data_o_50_), .Q_N(n1408), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_51_ (.CLK(clk), .D(n4077), .Q(data_o_51_), .Q_N(n1403), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_52_ (.CLK(clk), .D(n4076), .Q(data_o_52_), .Q_N(n1398), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_53_ (.CLK(clk), .D(n4075), .Q(data_o_53_), .Q_N(n1393), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_54_ (.CLK(clk), .D(n4074), .Q(data_o_54_), .Q_N(n1388), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_55_ (.CLK(clk), .D(n4073), .Q(data_o_55_), .Q_N(n1383), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_56_ (.CLK(clk), .D(n4072), .Q(data_o_56_), .Q_N(n1378), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_57_ (.CLK(clk), .D(n4071), .Q(data_o_57_), .Q_N(n1373), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_58_ (.CLK(clk), .D(n4070), .Q(data_o_58_), .Q_N(n1368), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_59_ (.CLK(clk), .D(n4069), .Q(data_o_59_), .Q_N(n1363), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_60_ (.CLK(clk), .D(n4068), .Q(data_o_60_), .Q_N(n1353), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_61_ (.CLK(clk), .D(n4067), .Q(data_o_61_), .Q_N(n1348), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_62_ (.CLK(clk), .D(n4066), .Q(data_o_62_), .Q_N(n1343), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_63_ (.CLK(clk), .D(n4065), .Q(data_o_63_), .Q_N(n1338), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_64_ (.CLK(clk), .D(n4064), .Q(data_o_64_), .Q_N(n1333), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_65_ (.CLK(clk), .D(n4063), .Q(data_o_65_), .Q_N(n1328), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_66_ (.CLK(clk), .D(n4062), .Q(data_o_66_), .Q_N(n1323), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_67_ (.CLK(clk), .D(n4061), .Q(data_o_67_), .Q_N(n1318), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_68_ (.CLK(clk), .D(n4060), .Q(data_o_68_), .Q_N(n1313), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_69_ (.CLK(clk), .D(n4059), .Q(data_o_69_), .Q_N(n1308), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_70_ (.CLK(clk), .D(n4058), .Q(data_o_70_), .Q_N(n1298), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_71_ (.CLK(clk), .D(n4057), .Q(data_o_71_), .Q_N(n1293), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_72_ (.CLK(clk), .D(n4056), .Q(data_o_72_), .Q_N(n1288), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_73_ (.CLK(clk), .D(n4055), .Q(data_o_73_), .Q_N(n1283), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_74_ (.CLK(clk), .D(n4054), .Q(data_o_74_), .Q_N(n1278), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_75_ (.CLK(clk), .D(n4053), .Q(data_o_75_), .Q_N(n1273), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_76_ (.CLK(clk), .D(n4052), .Q(data_o_76_), .Q_N(n1268), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_77_ (.CLK(clk), .D(n4051), .Q(data_o_77_), .Q_N(n1263), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_78_ (.CLK(clk), .D(n4050), .Q(data_o_78_), .Q_N(n1258), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_79_ (.CLK(clk), .D(n4049), .Q(data_o_79_), .Q_N(n1253), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_80_ (.CLK(clk), .D(n4048), .Q(data_o_80_), .Q_N(n1243), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_81_ (.CLK(clk), .D(n4047), .Q(data_o_81_), .Q_N(n1238), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_82_ (.CLK(clk), .D(n4046), .Q(data_o_82_), .Q_N(n1233), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_83_ (.CLK(clk), .D(n4045), .Q(data_o_83_), .Q_N(n1228), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_84_ (.CLK(clk), .D(n4044), .Q(data_o_84_), .Q_N(n1223), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_85_ (.CLK(clk), .D(n4043), .Q(data_o_85_), .Q_N(n1218), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_86_ (.CLK(clk), .D(n4042), .Q(data_o_86_), .Q_N(n1213), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_87_ (.CLK(clk), .D(n4041), .Q(data_o_87_), .Q_N(n1208), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_88_ (.CLK(clk), .D(n4040), .Q(data_o_88_), .Q_N(n1203), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_89_ (.CLK(clk), .D(n4039), .Q(data_o_89_), .Q_N(n1198), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_90_ (.CLK(clk), .D(n4038), .Q(data_o_90_), .Q_N(n1188), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_91_ (.CLK(clk), .D(n4037), .Q(data_o_91_), .Q_N(n1183), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_92_ (.CLK(clk), .D(n4036), .Q(data_o_92_), .Q_N(n1178), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_93_ (.CLK(clk), .D(n4035), .Q(data_o_93_), .Q_N(n1173), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_94_ (.CLK(clk), .D(n4034), .Q(data_o_94_), .Q_N(n1168), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_95_ (.CLK(clk), .D(n4033), .Q(data_o_95_), .Q_N(n1163), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_96_ (.CLK(clk), .D(n4032), .Q(data_o_96_), .Q_N(n1158), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_97_ (.CLK(clk), .D(n4031), .Q(data_o_97_), .Q_N(n1153), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_98_ (.CLK(clk), .D(n4030), .Q(data_o_98_), .Q_N(n1148), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_99_ (.CLK(clk), .D(n4028), .Q(data_o_99_), .Q_N(n1143), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_100_ (.CLK(clk), .D(n4027), .Q(data_o_100_), .Q_N(n1768), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_101_ (.CLK(clk), .D(n4026), .Q(data_o_101_), .Q_N(n1763), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_102_ (.CLK(clk), .D(n4025), .Q(data_o_102_), .Q_N(n1758), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_103_ (.CLK(clk), .D(n4024), .Q(data_o_103_), .Q_N(n1753), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_104_ (.CLK(clk), .D(n4023), .Q(data_o_104_), .Q_N(n1748), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_105_ (.CLK(clk), .D(n4022), .Q(data_o_105_), .Q_N(n1743), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_106_ (.CLK(clk), .D(n4021), .Q(data_o_106_), .Q_N(n1738), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_107_ (.CLK(clk), .D(n4020), .Q(data_o_107_), .Q_N(n1733), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_108_ (.CLK(clk), .D(n4019), .Q(data_o_108_), .Q_N(n1728), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_109_ (.CLK(clk), .D(n4018), .Q(data_o_109_), .Q_N(n1723), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_110_ (.CLK(clk), .D(n4017), .Q(data_o_110_), .Q_N(n1713), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_111_ (.CLK(clk), .D(n4016), .Q(data_o_111_), .Q_N(n1708), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_112_ (.CLK(clk), .D(n4015), .Q(data_o_112_), .Q_N(n1703), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_113_ (.CLK(clk), .D(n4014), .Q(data_o_113_), .Q_N(n1698), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_114_ (.CLK(clk), .D(n4013), .Q(data_o_114_), .Q_N(n1693), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_115_ (.CLK(clk), .D(n4012), .Q(data_o_115_), .Q_N(n1688), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_116_ (.CLK(clk), .D(n4011), .Q(data_o_116_), .Q_N(n1683), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_117_ (.CLK(clk), .D(n4010), .Q(data_o_117_), .Q_N(n1678), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_118_ (.CLK(clk), .D(n4009), .Q(data_o_118_), .Q_N(n1673), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_119_ (.CLK(clk), .D(n4008), .Q(data_o_119_), .Q_N(n1668), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_120_ (.CLK(clk), .D(n4007), .Q(data_o_120_), .Q_N(n1658), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_121_ (.CLK(clk), .D(n4006), .Q(data_o_121_), .Q_N(n1653), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_122_ (.CLK(clk), .D(n4005), .Q(data_o_122_), .Q_N(n1648), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_123_ (.CLK(clk), .D(n4004), .Q(data_o_123_), .Q_N(n1643), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_124_ (.CLK(clk), .D(n4003), .Q(data_o_124_), .Q_N(n1638), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_125_ (.CLK(clk), .D(n4002), .Q(data_o_125_), .Q_N(n1633), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_126_ (.CLK(clk), .D(n4001), .Q(data_o_126_), .Q_N(n1628), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_data_reg_reg_127_ (.CLK(clk), .D(n4134), .Q(data_o_127_), .Q_N(n1623), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_ready_o_reg (.CLK(clk), .D(next_addroundkey_ready_o), .Q(addroundkey_ready_o), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_round_reg_0_ (.CLK(clk), .D(n3938), .Q(addroundkey_round_0), .Q_N(n3736), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_round_reg_1_ (.CLK(clk), .D(n3937), .Q(addroundkey_round_1), .Q_N(net44327), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_round_reg_2_ (.CLK(clk), .D(n3936), .Q(addroundkey_round_2), .Q_N(net44332), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_round_reg_3_ (.CLK(clk), .D(n4136), .Q(addroundkey_round_3), .Q_N(net44340), .RESET_B(reset));
sg13g2_dfrbp_1 addroundkey_start_i_reg (.CLK(clk), .D(next_addroundkey_start_i), .Q(addroundkey_start_i), .RESET_B(reset));
sg13g2_dfrbp_2 first_round_reg_reg (.CLK(clk), .D(next_first_round_reg), .Q_N(n1115), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_0_ (.CLK(clk), .D(n4000), .Q(last_key_half_0), .Q_N(n3656), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_1_ (.CLK(clk), .D(n3999), .Q(last_key_half_1), .Q_N(n3654), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_2_ (.CLK(clk), .D(n3998), .Q(last_key_half_2), .Q_N(n3652), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_3_ (.CLK(clk), .D(n3997), .Q(last_key_half_3), .Q_N(n3650), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_4_ (.CLK(clk), .D(n3996), .Q(last_key_half_4), .Q_N(n3648), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_5_ (.CLK(clk), .D(n3995), .Q(last_key_half_5), .Q_N(n3646), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_6_ (.CLK(clk), .D(n3994), .Q(last_key_half_6), .Q_N(n3644), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_7_ (.CLK(clk), .D(n3993), .Q(last_key_half_7), .Q_N(n3642), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_8_ (.CLK(clk), .D(n3992), .Q(last_key_half_8), .Q_N(n3640), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_9_ (.CLK(clk), .D(n3991), .Q(last_key_half_9), .Q_N(n3638), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_10_ (.CLK(clk), .D(n3990), .Q(last_key_half_10), .Q_N(n3636), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_11_ (.CLK(clk), .D(n3989), .Q(last_key_half_11), .Q_N(n3634), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_12_ (.CLK(clk), .D(n3988), .Q(last_key_half_12), .Q_N(n3632), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_13_ (.CLK(clk), .D(n3987), .Q(last_key_half_13), .Q_N(n3630), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_14_ (.CLK(clk), .D(n3986), .Q(last_key_half_14), .Q_N(n3628), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_15_ (.CLK(clk), .D(n3985), .Q(last_key_half_15), .Q_N(n3626), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_16_ (.CLK(clk), .D(n3984), .Q(last_key_half_16), .Q_N(n3624), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_17_ (.CLK(clk), .D(n3983), .Q(last_key_half_17), .Q_N(n3622), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_18_ (.CLK(clk), .D(n3982), .Q(last_key_half_18), .Q_N(n3620), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_19_ (.CLK(clk), .D(n3981), .Q(last_key_half_19), .Q_N(n3618), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_20_ (.CLK(clk), .D(n3980), .Q(last_key_half_20), .Q_N(n3616), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_21_ (.CLK(clk), .D(n3979), .Q(last_key_half_21), .Q_N(n3614), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_22_ (.CLK(clk), .D(n3978), .Q(last_key_half_22), .Q_N(n3612), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_23_ (.CLK(clk), .D(n3977), .Q(last_key_half_23), .Q_N(n3610), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_24_ (.CLK(clk), .D(n3976), .Q(last_key_half_24), .Q_N(n3608), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_25_ (.CLK(clk), .D(n3975), .Q(last_key_half_25), .Q_N(n3606), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_26_ (.CLK(clk), .D(n3974), .Q(last_key_half_26), .Q_N(n3604), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_27_ (.CLK(clk), .D(n3973), .Q(last_key_half_27), .Q_N(n3602), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_28_ (.CLK(clk), .D(n3972), .Q(last_key_half_28), .Q_N(n3600), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_29_ (.CLK(clk), .D(n3971), .Q(last_key_half_29), .Q_N(n3598), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_30_ (.CLK(clk), .D(n3970), .Q(last_key_half_30), .Q_N(n3596), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_31_ (.CLK(clk), .D(n3969), .Q(last_key_half_31), .Q_N(n3594), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_32_ (.CLK(clk), .D(n3968), .Q(last_key_half_32), .Q_N(n3592), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_33_ (.CLK(clk), .D(n3967), .Q(last_key_half_33), .Q_N(n3590), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_34_ (.CLK(clk), .D(n3966), .Q(last_key_half_34), .Q_N(n3588), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_35_ (.CLK(clk), .D(n3965), .Q(last_key_half_35), .Q_N(n3586), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_36_ (.CLK(clk), .D(n3964), .Q(last_key_half_36), .Q_N(n3584), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_37_ (.CLK(clk), .D(n3963), .Q(last_key_half_37), .Q_N(n3582), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_38_ (.CLK(clk), .D(n3962), .Q(last_key_half_38), .Q_N(n3580), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_39_ (.CLK(clk), .D(n3961), .Q(last_key_half_39), .Q_N(n3578), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_40_ (.CLK(clk), .D(n3960), .Q(last_key_half_40), .Q_N(n3576), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_41_ (.CLK(clk), .D(n3959), .Q(last_key_half_41), .Q_N(n3574), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_42_ (.CLK(clk), .D(n3958), .Q(last_key_half_42), .Q_N(n3572), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_43_ (.CLK(clk), .D(n3957), .Q(last_key_half_43), .Q_N(n3570), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_44_ (.CLK(clk), .D(n3956), .Q(last_key_half_44), .Q_N(n3568), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_45_ (.CLK(clk), .D(n3955), .Q(last_key_half_45), .Q_N(n3566), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_46_ (.CLK(clk), .D(n3954), .Q(last_key_half_46), .Q_N(n3564), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_47_ (.CLK(clk), .D(n3953), .Q(last_key_half_47), .Q_N(n3562), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_48_ (.CLK(clk), .D(n3952), .Q(last_key_half_48), .Q_N(n3560), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_49_ (.CLK(clk), .D(n3951), .Q(last_key_half_49), .Q_N(n3558), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_50_ (.CLK(clk), .D(n3950), .Q(last_key_half_50), .Q_N(n3556), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_51_ (.CLK(clk), .D(n3949), .Q(last_key_half_51), .Q_N(n3554), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_52_ (.CLK(clk), .D(n3948), .Q(last_key_half_52), .Q_N(n3552), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_53_ (.CLK(clk), .D(n3947), .Q(last_key_half_53), .Q_N(n3550), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_54_ (.CLK(clk), .D(n3946), .Q(last_key_half_54), .Q_N(n3548), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_55_ (.CLK(clk), .D(n3945), .Q(last_key_half_55), .Q_N(n3546), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_56_ (.CLK(clk), .D(n3944), .Q(last_key_half_56), .Q_N(n3544), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_57_ (.CLK(clk), .D(n3943), .Q(last_key_half_57), .Q_N(n3542), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_58_ (.CLK(clk), .D(n3942), .Q(last_key_half_58), .Q_N(n3540), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_59_ (.CLK(clk), .D(n3941), .Q(last_key_half_59), .Q_N(n3538), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_60_ (.CLK(clk), .D(n3940), .Q(last_key_half_60), .Q_N(n3536), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_61_ (.CLK(clk), .D(n3939), .Q(last_key_half_61), .Q_N(n3534), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_62_ (.CLK(clk), .D(n4029), .Q(last_key_half_62), .Q_N(n3532), .RESET_B(reset));
sg13g2_dfrbp_1 last_key_half_reg_63_ (.CLK(clk), .D(n4135), .Q(last_key_half_63), .Q_N(n3530), .RESET_B(reset));
sg13g2_inv_4 r370_U23 (.A(r370_n21), .Y(r370_n19));
sg13g2_xnor2_1 r370_U25 (.A(r370_n26), .B(addroundkey_round_0), .Y(r370_n21));
sg13g2_xnor2_1 r371_U25 (.A(three_0), .B(addroundkey_round_0), .Y(r371_n21));
sg13g2_inv_4 r371_U23 (.A(r371_n21), .Y(r371_n19));
sg13g2_nor2_2 r371_U3 (.A(r371_n10), .B(r371_n12), .Y(N1323));
sg13g2_nor2_2 r372_U3 (.A(n4294), .B(r372_n12), .Y(N1324));
sg13g2_inv_4 r372_U23 (.A(r372_n21), .Y(r372_n19));
sg13g2_xnor2_1 r372_U25 (.A(r370_n26), .B(addroundkey_round_0), .Y(r372_n21));
sg13g2_nor2_2 r373_U3 (.A(r373_n12), .B(r373_n10), .Y(N1325));
sg13g2_xnor2_1 r373_U19 (.A(net26538), .B(addroundkey_round_2), .Y(r373_n15));
sg13g2_inv_4 r373_U31 (.A(net25972), .Y(r373_n26));
sg13g2_nand2_2 r373_U15 (.A(r373_n13), .B(r373_n19), .Y(r373_n12));
sg13g2_dfrbp_1 ready_o_reg (.CLK(clk), .D(next_ready_o), .Q(ready_o), .RESET_B(reset));
sg13g2_dfrbp_2 round_reg_0_ (.CLK(clk), .D(n4129), .Q(two_0), .Q_N(net47625), .RESET_B(reset));
sg13g2_dfrbp_1 round_reg_1_ (.CLK(clk), .D(n4130), .Q(four_1), .Q_N(net25927), .RESET_B(reset));
sg13g2_dfrbp_1 round_reg_2_ (.CLK(clk), .D(n4131), .Q(round_2_), .Q_N(net26537), .RESET_B(reset));
sg13g2_dfrbp_2 round_reg_3_ (.CLK(clk), .D(n4133), .Q_N(net47651), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg (.CLK(clk), .D(n4132), .Q(state), .Q_N(n4331), .RESET_B(reset));
keysched192 ks1(.clk(clk), .last_key_i_0_(keysched_last_key_i_0), .last_key_i_1_(keysched_last_key_i_1), .last_key_i_2_(keysched_last_key_i_2), .last_key_i_3_(keysched_last_key_i_3), .last_key_i_4_(keysched_last_key_i_4), .last_key_i_5_(keysched_last_key_i_5), .last_key_i_6_(keysched_last_key_i_6), .last_key_i_7_(keysched_last_key_i_7), .last_key_i_8_(keysched_last_key_i_8), .last_key_i_9_(keysched_last_key_i_9), .last_key_i_10_(keysched_last_key_i_10), .last_key_i_11_(keysched_last_key_i_11), .last_key_i_12_(keysched_last_key_i_12), .last_key_i_13_(keysched_last_key_i_13), .last_key_i_14_(keysched_last_key_i_14), .last_key_i_15_(keysched_last_key_i_15), .last_key_i_16_(keysched_last_key_i_16), .last_key_i_17_(keysched_last_key_i_17), .last_key_i_18_(keysched_last_key_i_18), .last_key_i_19_(keysched_last_key_i_19), .last_key_i_20_(keysched_last_key_i_20), .last_key_i_21_(keysched_last_key_i_21), .last_key_i_22_(keysched_last_key_i_22), .last_key_i_23_(keysched_last_key_i_23), .last_key_i_24_(keysched_last_key_i_24), .last_key_i_25_(keysched_last_key_i_25), .last_key_i_26_(keysched_last_key_i_26), .last_key_i_27_(keysched_last_key_i_27), .last_key_i_28_(keysched_last_key_i_28), .last_key_i_29_(keysched_last_key_i_29), .last_key_i_30_(keysched_last_key_i_30), .last_key_i_31_(keysched_last_key_i_31), .last_key_i_32_(keysched_last_key_i_32), .last_key_i_33_(keysched_last_key_i_33), .last_key_i_34_(keysched_last_key_i_34), .last_key_i_35_(keysched_last_key_i_35), .last_key_i_36_(keysched_last_key_i_36), .last_key_i_37_(keysched_last_key_i_37), .last_key_i_38_(keysched_last_key_i_38), .last_key_i_39_(keysched_last_key_i_39), .last_key_i_40_(keysched_last_key_i_40), .last_key_i_41_(keysched_last_key_i_41), .last_key_i_42_(keysched_last_key_i_42), .last_key_i_43_(keysched_last_key_i_43), .last_key_i_44_(keysched_last_key_i_44), .last_key_i_45_(keysched_last_key_i_45), .last_key_i_46_(keysched_last_key_i_46), .last_key_i_47_(keysched_last_key_i_47), .last_key_i_48_(keysched_last_key_i_48), .last_key_i_49_(keysched_last_key_i_49), .last_key_i_50_(keysched_last_key_i_50), .last_key_i_51_(keysched_last_key_i_51), .last_key_i_52_(keysched_last_key_i_52), .last_key_i_53_(keysched_last_key_i_53), .last_key_i_54_(keysched_last_key_i_54), .last_key_i_55_(keysched_last_key_i_55), .last_key_i_56_(keysched_last_key_i_56), .last_key_i_57_(keysched_last_key_i_57), .last_key_i_58_(keysched_last_key_i_58), .last_key_i_59_(keysched_last_key_i_59), .last_key_i_60_(keysched_last_key_i_60), .last_key_i_61_(keysched_last_key_i_61), .last_key_i_62_(keysched_last_key_i_62), .last_key_i_63_(keysched_last_key_i_63), .last_key_i_64_(keysched_last_key_i_64), .last_key_i_65_(keysched_last_key_i_65), .last_key_i_66_(keysched_last_key_i_66), .last_key_i_67_(keysched_last_key_i_67), .last_key_i_68_(keysched_last_key_i_68), .last_key_i_69_(keysched_last_key_i_69), .last_key_i_70_(keysched_last_key_i_70), .last_key_i_71_(keysched_last_key_i_71), .last_key_i_72_(keysched_last_key_i_72), .last_key_i_73_(keysched_last_key_i_73), .last_key_i_74_(keysched_last_key_i_74), .last_key_i_75_(keysched_last_key_i_75), .last_key_i_76_(keysched_last_key_i_76), .last_key_i_77_(keysched_last_key_i_77), .last_key_i_78_(keysched_last_key_i_78), .last_key_i_79_(keysched_last_key_i_79), .last_key_i_80_(keysched_last_key_i_80), .last_key_i_81_(keysched_last_key_i_81), .last_key_i_82_(keysched_last_key_i_82), .last_key_i_83_(keysched_last_key_i_83), .last_key_i_84_(keysched_last_key_i_84), .last_key_i_85_(keysched_last_key_i_85), .last_key_i_86_(keysched_last_key_i_86), .last_key_i_87_(keysched_last_key_i_87), .last_key_i_88_(keysched_last_key_i_88), .last_key_i_89_(keysched_last_key_i_89), .last_key_i_90_(keysched_last_key_i_90), .last_key_i_91_(keysched_last_key_i_91), .last_key_i_92_(keysched_last_key_i_92), .last_key_i_93_(keysched_last_key_i_93), .last_key_i_94_(keysched_last_key_i_94), .last_key_i_95_(keysched_last_key_i_95), .last_key_i_96_(keysched_last_key_i_96), .last_key_i_97_(keysched_last_key_i_97), .last_key_i_98_(keysched_last_key_i_98), .last_key_i_99_(keysched_last_key_i_99), .last_key_i_100_(keysched_last_key_i_100), .last_key_i_101_(keysched_last_key_i_101), .last_key_i_102_(keysched_last_key_i_102), .last_key_i_103_(keysched_last_key_i_103), .last_key_i_104_(keysched_last_key_i_104), .last_key_i_105_(keysched_last_key_i_105), .last_key_i_106_(keysched_last_key_i_106), .last_key_i_107_(keysched_last_key_i_107), .last_key_i_108_(keysched_last_key_i_108), .last_key_i_109_(keysched_last_key_i_109), .last_key_i_110_(keysched_last_key_i_110), .last_key_i_111_(keysched_last_key_i_111), .last_key_i_112_(keysched_last_key_i_112), .last_key_i_113_(keysched_last_key_i_113), .last_key_i_114_(keysched_last_key_i_114), .last_key_i_115_(keysched_last_key_i_115), .last_key_i_116_(keysched_last_key_i_116), .last_key_i_117_(keysched_last_key_i_117), .last_key_i_118_(keysched_last_key_i_118), .last_key_i_119_(keysched_last_key_i_119), .last_key_i_120_(keysched_last_key_i_120), .last_key_i_121_(keysched_last_key_i_121), .last_key_i_122_(keysched_last_key_i_122), .last_key_i_123_(keysched_last_key_i_123), .last_key_i_124_(keysched_last_key_i_124), .last_key_i_125_(keysched_last_key_i_125), .last_key_i_126_(keysched_last_key_i_126), .last_key_i_127_(keysched_last_key_i_127), .last_key_i_128_(keysched_last_key_i_128), .last_key_i_129_(keysched_last_key_i_129), .last_key_i_130_(keysched_last_key_i_130), .last_key_i_131_(keysched_last_key_i_131), .last_key_i_132_(keysched_last_key_i_132), .last_key_i_133_(keysched_last_key_i_133), .last_key_i_134_(keysched_last_key_i_134), .last_key_i_135_(keysched_last_key_i_135), .last_key_i_136_(keysched_last_key_i_136), .last_key_i_137_(keysched_last_key_i_137), .last_key_i_138_(keysched_last_key_i_138), .last_key_i_139_(keysched_last_key_i_139), .last_key_i_140_(keysched_last_key_i_140), .last_key_i_141_(keysched_last_key_i_141), .last_key_i_142_(keysched_last_key_i_142), .last_key_i_143_(keysched_last_key_i_143), .last_key_i_144_(keysched_last_key_i_144), .last_key_i_145_(keysched_last_key_i_145), .last_key_i_146_(keysched_last_key_i_146), .last_key_i_147_(keysched_last_key_i_147), .last_key_i_148_(keysched_last_key_i_148), .last_key_i_149_(keysched_last_key_i_149), .last_key_i_150_(keysched_last_key_i_150), .last_key_i_151_(keysched_last_key_i_151), .last_key_i_152_(keysched_last_key_i_152), .last_key_i_153_(keysched_last_key_i_153), .last_key_i_154_(keysched_last_key_i_154), .last_key_i_155_(keysched_last_key_i_155), .last_key_i_156_(keysched_last_key_i_156), .last_key_i_157_(keysched_last_key_i_157), .last_key_i_158_(keysched_last_key_i_158), .last_key_i_159_(keysched_last_key_i_159), .last_key_i_160_(keysched_last_key_i_160), .last_key_i_161_(keysched_last_key_i_161), .last_key_i_162_(keysched_last_key_i_162), .last_key_i_163_(keysched_last_key_i_163), .last_key_i_164_(keysched_last_key_i_164), .last_key_i_165_(keysched_last_key_i_165), .last_key_i_166_(keysched_last_key_i_166), .last_key_i_167_(keysched_last_key_i_167), .last_key_i_168_(keysched_last_key_i_168), .last_key_i_169_(keysched_last_key_i_169), .last_key_i_170_(keysched_last_key_i_170), .last_key_i_171_(keysched_last_key_i_171), .last_key_i_172_(keysched_last_key_i_172), .last_key_i_173_(keysched_last_key_i_173), .last_key_i_174_(keysched_last_key_i_174), .last_key_i_175_(keysched_last_key_i_175), .last_key_i_176_(keysched_last_key_i_176), .last_key_i_177_(keysched_last_key_i_177), .last_key_i_178_(keysched_last_key_i_178), .last_key_i_179_(keysched_last_key_i_179), .last_key_i_180_(keysched_last_key_i_180), .last_key_i_181_(keysched_last_key_i_181), .last_key_i_182_(keysched_last_key_i_182), .last_key_i_183_(keysched_last_key_i_183), .last_key_i_184_(keysched_last_key_i_184), .last_key_i_185_(keysched_last_key_i_185), .last_key_i_186_(keysched_last_key_i_186), .last_key_i_187_(keysched_last_key_i_187), .last_key_i_188_(keysched_last_key_i_188), .last_key_i_189_(keysched_last_key_i_189), .last_key_i_190_(keysched_last_key_i_190), .last_key_i_191_(keysched_last_key_i_191), .new_key_o_0_(keysched_new_key_o_0), .new_key_o_1_(keysched_new_key_o_1), .new_key_o_2_(keysched_new_key_o_2), .new_key_o_3_(keysched_new_key_o_3), .new_key_o_4_(keysched_new_key_o_4), .new_key_o_5_(keysched_new_key_o_5), .new_key_o_6_(keysched_new_key_o_6), .new_key_o_7_(keysched_new_key_o_7), .new_key_o_8_(keysched_new_key_o_8), .new_key_o_9_(keysched_new_key_o_9), .new_key_o_10_(keysched_new_key_o_10), .new_key_o_11_(keysched_new_key_o_11), .new_key_o_12_(keysched_new_key_o_12), .new_key_o_13_(keysched_new_key_o_13), .new_key_o_14_(keysched_new_key_o_14), .new_key_o_15_(keysched_new_key_o_15), .new_key_o_16_(keysched_new_key_o_16), .new_key_o_17_(keysched_new_key_o_17), .new_key_o_18_(keysched_new_key_o_18), .new_key_o_19_(keysched_new_key_o_19), .new_key_o_20_(keysched_new_key_o_20), .new_key_o_21_(keysched_new_key_o_21), .new_key_o_22_(keysched_new_key_o_22), .new_key_o_23_(keysched_new_key_o_23), .new_key_o_24_(keysched_new_key_o_24), .new_key_o_25_(keysched_new_key_o_25), .new_key_o_26_(keysched_new_key_o_26), .new_key_o_27_(keysched_new_key_o_27), .new_key_o_28_(keysched_new_key_o_28), .new_key_o_29_(keysched_new_key_o_29), .new_key_o_30_(keysched_new_key_o_30), .new_key_o_31_(keysched_new_key_o_31), .new_key_o_32_(keysched_new_key_o_32), .new_key_o_33_(keysched_new_key_o_33), .new_key_o_34_(keysched_new_key_o_34), .new_key_o_35_(keysched_new_key_o_35), .new_key_o_36_(keysched_new_key_o_36), .new_key_o_37_(keysched_new_key_o_37), .new_key_o_38_(keysched_new_key_o_38), .new_key_o_39_(keysched_new_key_o_39), .new_key_o_40_(keysched_new_key_o_40), .new_key_o_41_(keysched_new_key_o_41), .new_key_o_42_(keysched_new_key_o_42), .new_key_o_43_(keysched_new_key_o_43), .new_key_o_44_(keysched_new_key_o_44), .new_key_o_45_(keysched_new_key_o_45), .new_key_o_46_(keysched_new_key_o_46), .new_key_o_47_(keysched_new_key_o_47), .new_key_o_48_(keysched_new_key_o_48), .new_key_o_49_(keysched_new_key_o_49), .new_key_o_50_(keysched_new_key_o_50), .new_key_o_51_(keysched_new_key_o_51), .new_key_o_52_(keysched_new_key_o_52), .new_key_o_53_(keysched_new_key_o_53), .new_key_o_54_(keysched_new_key_o_54), .new_key_o_55_(keysched_new_key_o_55), .new_key_o_56_(keysched_new_key_o_56), .new_key_o_57_(keysched_new_key_o_57), .new_key_o_58_(keysched_new_key_o_58), .new_key_o_59_(keysched_new_key_o_59), .new_key_o_60_(keysched_new_key_o_60), .new_key_o_61_(keysched_new_key_o_61), .new_key_o_62_(keysched_new_key_o_62), .new_key_o_63_(keysched_new_key_o_63), .new_key_o_64_(keysched_new_key_o_64), .new_key_o_65_(keysched_new_key_o_65), .new_key_o_66_(keysched_new_key_o_66), .new_key_o_67_(keysched_new_key_o_67), .new_key_o_68_(keysched_new_key_o_68), .new_key_o_69_(keysched_new_key_o_69), .new_key_o_70_(keysched_new_key_o_70), .new_key_o_71_(keysched_new_key_o_71), .new_key_o_72_(keysched_new_key_o_72), .new_key_o_73_(keysched_new_key_o_73), .new_key_o_74_(keysched_new_key_o_74), .new_key_o_75_(keysched_new_key_o_75), .new_key_o_76_(keysched_new_key_o_76), .new_key_o_77_(keysched_new_key_o_77), .new_key_o_78_(keysched_new_key_o_78), .new_key_o_79_(keysched_new_key_o_79), .new_key_o_80_(keysched_new_key_o_80), .new_key_o_81_(keysched_new_key_o_81), .new_key_o_82_(keysched_new_key_o_82), .new_key_o_83_(keysched_new_key_o_83), .new_key_o_84_(keysched_new_key_o_84), .new_key_o_85_(keysched_new_key_o_85), .new_key_o_86_(keysched_new_key_o_86), .new_key_o_87_(keysched_new_key_o_87), .new_key_o_88_(keysched_new_key_o_88), .new_key_o_89_(keysched_new_key_o_89), .new_key_o_90_(keysched_new_key_o_90), .new_key_o_91_(keysched_new_key_o_91), .new_key_o_92_(keysched_new_key_o_92), .new_key_o_93_(keysched_new_key_o_93), .new_key_o_94_(keysched_new_key_o_94), .new_key_o_95_(keysched_new_key_o_95), .new_key_o_96_(keysched_new_key_o_96), .new_key_o_97_(keysched_new_key_o_97), .new_key_o_98_(keysched_new_key_o_98), .new_key_o_99_(keysched_new_key_o_99), .new_key_o_100_(keysched_new_key_o_100), .new_key_o_101_(keysched_new_key_o_101), .new_key_o_102_(keysched_new_key_o_102), .new_key_o_103_(keysched_new_key_o_103), .new_key_o_104_(keysched_new_key_o_104), .new_key_o_105_(keysched_new_key_o_105), .new_key_o_106_(keysched_new_key_o_106), .new_key_o_107_(keysched_new_key_o_107), .new_key_o_108_(keysched_new_key_o_108), .new_key_o_109_(keysched_new_key_o_109), .new_key_o_110_(keysched_new_key_o_110), .new_key_o_111_(keysched_new_key_o_111), .new_key_o_112_(keysched_new_key_o_112), .new_key_o_113_(keysched_new_key_o_113), .new_key_o_114_(keysched_new_key_o_114), .new_key_o_115_(keysched_new_key_o_115), .new_key_o_116_(keysched_new_key_o_116), .new_key_o_117_(keysched_new_key_o_117), .new_key_o_118_(keysched_new_key_o_118), .new_key_o_119_(keysched_new_key_o_119), .new_key_o_120_(keysched_new_key_o_120), .new_key_o_121_(keysched_new_key_o_121), .new_key_o_122_(keysched_new_key_o_122), .new_key_o_123_(keysched_new_key_o_123), .new_key_o_124_(keysched_new_key_o_124), .new_key_o_125_(keysched_new_key_o_125), .new_key_o_126_(keysched_new_key_o_126), .new_key_o_127_(keysched_new_key_o_127), .new_key_o_128_(keysched_new_key_o_128), .new_key_o_129_(keysched_new_key_o_129), .new_key_o_130_(keysched_new_key_o_130), .new_key_o_131_(keysched_new_key_o_131), .new_key_o_132_(keysched_new_key_o_132), .new_key_o_133_(keysched_new_key_o_133), .new_key_o_134_(keysched_new_key_o_134), .new_key_o_135_(keysched_new_key_o_135), .new_key_o_136_(keysched_new_key_o_136), .new_key_o_137_(keysched_new_key_o_137), .new_key_o_138_(keysched_new_key_o_138), .new_key_o_139_(keysched_new_key_o_139), .new_key_o_140_(keysched_new_key_o_140), .new_key_o_141_(keysched_new_key_o_141), .new_key_o_142_(keysched_new_key_o_142), .new_key_o_143_(keysched_new_key_o_143), .new_key_o_144_(keysched_new_key_o_144), .new_key_o_145_(keysched_new_key_o_145), .new_key_o_146_(keysched_new_key_o_146), .new_key_o_147_(keysched_new_key_o_147), .new_key_o_148_(keysched_new_key_o_148), .new_key_o_149_(keysched_new_key_o_149), .new_key_o_150_(keysched_new_key_o_150), .new_key_o_151_(keysched_new_key_o_151), .new_key_o_152_(keysched_new_key_o_152), .new_key_o_153_(keysched_new_key_o_153), .new_key_o_154_(keysched_new_key_o_154), .new_key_o_155_(keysched_new_key_o_155), .new_key_o_156_(keysched_new_key_o_156), .new_key_o_157_(keysched_new_key_o_157), .new_key_o_158_(keysched_new_key_o_158), .new_key_o_159_(keysched_new_key_o_159), .new_key_o_160_(keysched_new_key_o_160), .new_key_o_161_(keysched_new_key_o_161), .new_key_o_162_(keysched_new_key_o_162), .new_key_o_163_(keysched_new_key_o_163), .new_key_o_164_(keysched_new_key_o_164), .new_key_o_165_(keysched_new_key_o_165), .new_key_o_166_(keysched_new_key_o_166), .new_key_o_167_(keysched_new_key_o_167), .new_key_o_168_(keysched_new_key_o_168), .new_key_o_169_(keysched_new_key_o_169), .new_key_o_170_(keysched_new_key_o_170), .new_key_o_171_(keysched_new_key_o_171), .new_key_o_172_(keysched_new_key_o_172), .new_key_o_173_(keysched_new_key_o_173), .new_key_o_174_(keysched_new_key_o_174), .new_key_o_175_(keysched_new_key_o_175), .new_key_o_176_(keysched_new_key_o_176), .new_key_o_177_(keysched_new_key_o_177), .new_key_o_178_(keysched_new_key_o_178), .new_key_o_179_(keysched_new_key_o_179), .new_key_o_180_(keysched_new_key_o_180), .new_key_o_181_(keysched_new_key_o_181), .new_key_o_182_(keysched_new_key_o_182), .new_key_o_183_(keysched_new_key_o_183), .new_key_o_184_(keysched_new_key_o_184), .new_key_o_185_(keysched_new_key_o_185), .new_key_o_186_(keysched_new_key_o_186), .new_key_o_187_(keysched_new_key_o_187), .new_key_o_188_(keysched_new_key_o_188), .new_key_o_189_(keysched_new_key_o_189), .new_key_o_190_(keysched_new_key_o_190), .new_key_o_191_(keysched_new_key_o_191), .ready_o(keysched_ready_o), .reset(reset), .round_i_0_(keysched_round_i_0), .round_i_1_(keysched_round_i_1), .round_i_2_(keysched_round_i_2), .round_i_3_(keysched_round_i_3), .sbox_access_o(keysched_sbox_access_o), .sbox_data_i_0_(n4276), .sbox_data_i_1_(sbox_data_o_1), .sbox_data_i_2_(sbox_data_o_2), .sbox_data_i_3_(n4289), .sbox_data_i_4_(sbox_data_o_4), .sbox_data_i_5_(sbox_data_o_5), .sbox_data_i_6_(sbox_data_o_6), .sbox_data_i_7_(sbox_data_o_7), .sbox_data_o_0_(keysched_sbox_data_o_0), .sbox_data_o_1_(keysched_sbox_data_o_1), .sbox_data_o_2_(keysched_sbox_data_o_2), .sbox_data_o_3_(keysched_sbox_data_o_3), .sbox_data_o_4_(keysched_sbox_data_o_4), .sbox_data_o_5_(keysched_sbox_data_o_5), .sbox_data_o_6_(keysched_sbox_data_o_6), .sbox_data_o_7_(keysched_sbox_data_o_7), .sbox_decrypt_o(), .start_i(keysched_start_i));
mixcolum mix1(.clk(clk), .data_i_0_(mixcol_data_i_0), .data_i_1_(mixcol_data_i_1), .data_i_2_(mixcol_data_i_2), .data_i_3_(mixcol_data_i_3), .data_i_4_(mixcol_data_i_4), .data_i_5_(mixcol_data_i_5), .data_i_6_(mixcol_data_i_6), .data_i_7_(mixcol_data_i_7), .data_i_8_(mixcol_data_i_8), .data_i_9_(mixcol_data_i_9), .data_i_10_(mixcol_data_i_10), .data_i_11_(mixcol_data_i_11), .data_i_12_(mixcol_data_i_12), .data_i_13_(mixcol_data_i_13), .data_i_14_(mixcol_data_i_14), .data_i_15_(mixcol_data_i_15), .data_i_16_(mixcol_data_i_16), .data_i_17_(mixcol_data_i_17), .data_i_18_(mixcol_data_i_18), .data_i_19_(mixcol_data_i_19), .data_i_20_(mixcol_data_i_20), .data_i_21_(mixcol_data_i_21), .data_i_22_(mixcol_data_i_22), .data_i_23_(mixcol_data_i_23), .data_i_24_(mixcol_data_i_24), .data_i_25_(mixcol_data_i_25), .data_i_26_(mixcol_data_i_26), .data_i_27_(mixcol_data_i_27), .data_i_28_(mixcol_data_i_28), .data_i_29_(mixcol_data_i_29), .data_i_30_(mixcol_data_i_30), .data_i_31_(mixcol_data_i_31), .data_i_32_(mixcol_data_i_32), .data_i_33_(mixcol_data_i_33), .data_i_34_(mixcol_data_i_34), .data_i_35_(mixcol_data_i_35), .data_i_36_(mixcol_data_i_36), .data_i_37_(mixcol_data_i_37), .data_i_38_(mixcol_data_i_38), .data_i_39_(mixcol_data_i_39), .data_i_40_(mixcol_data_i_40), .data_i_41_(mixcol_data_i_41), .data_i_42_(mixcol_data_i_42), .data_i_43_(mixcol_data_i_43), .data_i_44_(mixcol_data_i_44), .data_i_45_(mixcol_data_i_45), .data_i_46_(mixcol_data_i_46), .data_i_47_(mixcol_data_i_47), .data_i_48_(mixcol_data_i_48), .data_i_49_(mixcol_data_i_49), .data_i_50_(mixcol_data_i_50), .data_i_51_(mixcol_data_i_51), .data_i_52_(mixcol_data_i_52), .data_i_53_(mixcol_data_i_53), .data_i_54_(mixcol_data_i_54), .data_i_55_(mixcol_data_i_55), .data_i_56_(mixcol_data_i_56), .data_i_57_(mixcol_data_i_57), .data_i_58_(mixcol_data_i_58), .data_i_59_(mixcol_data_i_59), .data_i_60_(mixcol_data_i_60), .data_i_61_(mixcol_data_i_61), .data_i_62_(mixcol_data_i_62), .data_i_63_(mixcol_data_i_63), .data_i_64_(mixcol_data_i_64), .data_i_65_(mixcol_data_i_65), .data_i_66_(mixcol_data_i_66), .data_i_67_(mixcol_data_i_67), .data_i_68_(mixcol_data_i_68), .data_i_69_(mixcol_data_i_69), .data_i_70_(mixcol_data_i_70), .data_i_71_(mixcol_data_i_71), .data_i_72_(mixcol_data_i_72), .data_i_73_(mixcol_data_i_73), .data_i_74_(mixcol_data_i_74), .data_i_75_(mixcol_data_i_75), .data_i_76_(mixcol_data_i_76), .data_i_77_(mixcol_data_i_77), .data_i_78_(mixcol_data_i_78), .data_i_79_(mixcol_data_i_79), .data_i_80_(mixcol_data_i_80), .data_i_81_(mixcol_data_i_81), .data_i_82_(mixcol_data_i_82), .data_i_83_(mixcol_data_i_83), .data_i_84_(mixcol_data_i_84), .data_i_85_(mixcol_data_i_85), .data_i_86_(mixcol_data_i_86), .data_i_87_(mixcol_data_i_87), .data_i_88_(mixcol_data_i_88), .data_i_89_(mixcol_data_i_89), .data_i_90_(mixcol_data_i_90), .data_i_91_(mixcol_data_i_91), .data_i_92_(mixcol_data_i_92), .data_i_93_(mixcol_data_i_93), .data_i_94_(mixcol_data_i_94), .data_i_95_(mixcol_data_i_95), .data_i_96_(mixcol_data_i_96), .data_i_97_(mixcol_data_i_97), .data_i_98_(mixcol_data_i_98), .data_i_99_(mixcol_data_i_99), .data_i_100_(mixcol_data_i_100), .data_i_101_(mixcol_data_i_101), .data_i_102_(mixcol_data_i_102), .data_i_103_(mixcol_data_i_103), .data_i_104_(mixcol_data_i_104), .data_i_105_(mixcol_data_i_105), .data_i_106_(mixcol_data_i_106), .data_i_107_(mixcol_data_i_107), .data_i_108_(mixcol_data_i_108), .data_i_109_(mixcol_data_i_109), .data_i_110_(mixcol_data_i_110), .data_i_111_(mixcol_data_i_111), .data_i_112_(mixcol_data_i_112), .data_i_113_(mixcol_data_i_113), .data_i_114_(mixcol_data_i_114), .data_i_115_(mixcol_data_i_115), .data_i_116_(mixcol_data_i_116), .data_i_117_(mixcol_data_i_117), .data_i_118_(mixcol_data_i_118), .data_i_119_(mixcol_data_i_119), .data_i_120_(mixcol_data_i_120), .data_i_121_(mixcol_data_i_121), .data_i_122_(mixcol_data_i_122), .data_i_123_(mixcol_data_i_123), .data_i_124_(mixcol_data_i_124), .data_i_125_(mixcol_data_i_125), .data_i_126_(mixcol_data_i_126), .data_i_127_(mixcol_data_i_127), .data_o_0_(mixcol_data_o_0), .data_o_1_(mixcol_data_o_1), .data_o_2_(mixcol_data_o_2), .data_o_3_(mixcol_data_o_3), .data_o_4_(mixcol_data_o_4), .data_o_5_(mixcol_data_o_5), .data_o_6_(mixcol_data_o_6), .data_o_7_(mixcol_data_o_7), .data_o_8_(mixcol_data_o_8), .data_o_9_(mixcol_data_o_9), .data_o_10_(mixcol_data_o_10), .data_o_11_(mixcol_data_o_11), .data_o_12_(mixcol_data_o_12), .data_o_13_(mixcol_data_o_13), .data_o_14_(mixcol_data_o_14), .data_o_15_(mixcol_data_o_15), .data_o_16_(mixcol_data_o_16), .data_o_17_(mixcol_data_o_17), .data_o_18_(mixcol_data_o_18), .data_o_19_(mixcol_data_o_19), .data_o_20_(mixcol_data_o_20), .data_o_21_(mixcol_data_o_21), .data_o_22_(mixcol_data_o_22), .data_o_23_(mixcol_data_o_23), .data_o_24_(mixcol_data_o_24), .data_o_25_(mixcol_data_o_25), .data_o_26_(mixcol_data_o_26), .data_o_27_(mixcol_data_o_27), .data_o_28_(mixcol_data_o_28), .data_o_29_(mixcol_data_o_29), .data_o_30_(mixcol_data_o_30), .data_o_31_(mixcol_data_o_31), .data_o_32_(mixcol_data_o_32), .data_o_33_(mixcol_data_o_33), .data_o_34_(mixcol_data_o_34), .data_o_35_(mixcol_data_o_35), .data_o_36_(mixcol_data_o_36), .data_o_37_(mixcol_data_o_37), .data_o_38_(mixcol_data_o_38), .data_o_39_(mixcol_data_o_39), .data_o_40_(mixcol_data_o_40), .data_o_41_(mixcol_data_o_41), .data_o_42_(mixcol_data_o_42), .data_o_43_(mixcol_data_o_43), .data_o_44_(mixcol_data_o_44), .data_o_45_(mixcol_data_o_45), .data_o_46_(mixcol_data_o_46), .data_o_47_(mixcol_data_o_47), .data_o_48_(mixcol_data_o_48), .data_o_49_(mixcol_data_o_49), .data_o_50_(mixcol_data_o_50), .data_o_51_(mixcol_data_o_51), .data_o_52_(mixcol_data_o_52), .data_o_53_(mixcol_data_o_53), .data_o_54_(mixcol_data_o_54), .data_o_55_(mixcol_data_o_55), .data_o_56_(mixcol_data_o_56), .data_o_57_(mixcol_data_o_57), .data_o_58_(mixcol_data_o_58), .data_o_59_(mixcol_data_o_59), .data_o_60_(mixcol_data_o_60), .data_o_61_(mixcol_data_o_61), .data_o_62_(mixcol_data_o_62), .data_o_63_(mixcol_data_o_63), .data_o_64_(mixcol_data_o_64), .data_o_65_(mixcol_data_o_65), .data_o_66_(mixcol_data_o_66), .data_o_67_(mixcol_data_o_67), .data_o_68_(mixcol_data_o_68), .data_o_69_(mixcol_data_o_69), .data_o_70_(mixcol_data_o_70), .data_o_71_(mixcol_data_o_71), .data_o_72_(mixcol_data_o_72), .data_o_73_(mixcol_data_o_73), .data_o_74_(mixcol_data_o_74), .data_o_75_(mixcol_data_o_75), .data_o_76_(mixcol_data_o_76), .data_o_77_(mixcol_data_o_77), .data_o_78_(mixcol_data_o_78), .data_o_79_(mixcol_data_o_79), .data_o_80_(mixcol_data_o_80), .data_o_81_(mixcol_data_o_81), .data_o_82_(mixcol_data_o_82), .data_o_83_(mixcol_data_o_83), .data_o_84_(mixcol_data_o_84), .data_o_85_(mixcol_data_o_85), .data_o_86_(mixcol_data_o_86), .data_o_87_(mixcol_data_o_87), .data_o_88_(mixcol_data_o_88), .data_o_89_(mixcol_data_o_89), .data_o_90_(mixcol_data_o_90), .data_o_91_(mixcol_data_o_91), .data_o_92_(mixcol_data_o_92), .data_o_93_(mixcol_data_o_93), .data_o_94_(mixcol_data_o_94), .data_o_95_(mixcol_data_o_95), .data_o_96_(mixcol_data_o_96), .data_o_97_(mixcol_data_o_97), .data_o_98_(mixcol_data_o_98), .data_o_99_(mixcol_data_o_99), .data_o_100_(mixcol_data_o_100), .data_o_101_(mixcol_data_o_101), .data_o_102_(mixcol_data_o_102), .data_o_103_(mixcol_data_o_103), .data_o_104_(mixcol_data_o_104), .data_o_105_(mixcol_data_o_105), .data_o_106_(mixcol_data_o_106), .data_o_107_(mixcol_data_o_107), .data_o_108_(mixcol_data_o_108), .data_o_109_(mixcol_data_o_109), .data_o_110_(mixcol_data_o_110), .data_o_111_(mixcol_data_o_111), .data_o_112_(mixcol_data_o_112), .data_o_113_(mixcol_data_o_113), .data_o_114_(mixcol_data_o_114), .data_o_115_(mixcol_data_o_115), .data_o_116_(mixcol_data_o_116), .data_o_117_(mixcol_data_o_117), .data_o_118_(mixcol_data_o_118), .data_o_119_(mixcol_data_o_119), .data_o_120_(mixcol_data_o_120), .data_o_121_(mixcol_data_o_121), .data_o_122_(mixcol_data_o_122), .data_o_123_(mixcol_data_o_123), .data_o_124_(mixcol_data_o_124), .data_o_125_(mixcol_data_o_125), .data_o_126_(mixcol_data_o_126), .data_o_127_(mixcol_data_o_127), .decrypt_i(decrypt_i), .ready_o(mixcol_ready_o), .reset(reset), .start_i(mixcol_start_i));
sbox sbox1(.clk(clk), .data_i_0_(sbox_data_i_0), .data_i_1_(sbox_data_i_1), .data_i_2_(sbox_data_i_2), .data_i_3_(sbox_data_i_3), .data_i_4_(sbox_data_i_4), .data_i_5_(sbox_data_i_5), .data_i_6_(sbox_data_i_6), .data_i_7_(sbox_data_i_7), .data_o_0_(sbox_data_o_0), .data_o_1_(sbox_data_o_1), .data_o_2_(sbox_data_o_2), .data_o_3_(sbox_data_o_3), .data_o_4_(sbox_data_o_4), .data_o_5_(sbox_data_o_5), .data_o_6_(sbox_data_o_6), .data_o_7_(sbox_data_o_7), .decrypt_i(sbox_decrypt_i), .reset(reset));
subbytes sub1(.clk(clk), .data_i_0_(subbytes_data_i_0), .data_i_1_(subbytes_data_i_1), .data_i_2_(subbytes_data_i_2), .data_i_3_(subbytes_data_i_3), .data_i_4_(subbytes_data_i_4), .data_i_5_(subbytes_data_i_5), .data_i_6_(subbytes_data_i_6), .data_i_7_(subbytes_data_i_7), .data_i_8_(subbytes_data_i_8), .data_i_9_(subbytes_data_i_9), .data_i_10_(subbytes_data_i_10), .data_i_11_(subbytes_data_i_11), .data_i_12_(subbytes_data_i_12), .data_i_13_(subbytes_data_i_13), .data_i_14_(subbytes_data_i_14), .data_i_15_(subbytes_data_i_15), .data_i_16_(subbytes_data_i_16), .data_i_17_(subbytes_data_i_17), .data_i_18_(subbytes_data_i_18), .data_i_19_(subbytes_data_i_19), .data_i_20_(subbytes_data_i_20), .data_i_21_(subbytes_data_i_21), .data_i_22_(subbytes_data_i_22), .data_i_23_(subbytes_data_i_23), .data_i_24_(subbytes_data_i_24), .data_i_25_(subbytes_data_i_25), .data_i_26_(subbytes_data_i_26), .data_i_27_(subbytes_data_i_27), .data_i_28_(subbytes_data_i_28), .data_i_29_(subbytes_data_i_29), .data_i_30_(subbytes_data_i_30), .data_i_31_(subbytes_data_i_31), .data_i_32_(subbytes_data_i_32), .data_i_33_(subbytes_data_i_33), .data_i_34_(subbytes_data_i_34), .data_i_35_(subbytes_data_i_35), .data_i_36_(subbytes_data_i_36), .data_i_37_(subbytes_data_i_37), .data_i_38_(subbytes_data_i_38), .data_i_39_(subbytes_data_i_39), .data_i_40_(subbytes_data_i_40), .data_i_41_(subbytes_data_i_41), .data_i_42_(subbytes_data_i_42), .data_i_43_(subbytes_data_i_43), .data_i_44_(subbytes_data_i_44), .data_i_45_(subbytes_data_i_45), .data_i_46_(subbytes_data_i_46), .data_i_47_(subbytes_data_i_47), .data_i_48_(subbytes_data_i_48), .data_i_49_(subbytes_data_i_49), .data_i_50_(subbytes_data_i_50), .data_i_51_(subbytes_data_i_51), .data_i_52_(subbytes_data_i_52), .data_i_53_(subbytes_data_i_53), .data_i_54_(subbytes_data_i_54), .data_i_55_(subbytes_data_i_55), .data_i_56_(subbytes_data_i_56), .data_i_57_(subbytes_data_i_57), .data_i_58_(subbytes_data_i_58), .data_i_59_(subbytes_data_i_59), .data_i_60_(subbytes_data_i_60), .data_i_61_(subbytes_data_i_61), .data_i_62_(subbytes_data_i_62), .data_i_63_(subbytes_data_i_63), .data_i_64_(subbytes_data_i_64), .data_i_65_(subbytes_data_i_65), .data_i_66_(subbytes_data_i_66), .data_i_67_(subbytes_data_i_67), .data_i_68_(subbytes_data_i_68), .data_i_69_(subbytes_data_i_69), .data_i_70_(subbytes_data_i_70), .data_i_71_(subbytes_data_i_71), .data_i_72_(subbytes_data_i_72), .data_i_73_(subbytes_data_i_73), .data_i_74_(subbytes_data_i_74), .data_i_75_(subbytes_data_i_75), .data_i_76_(subbytes_data_i_76), .data_i_77_(subbytes_data_i_77), .data_i_78_(subbytes_data_i_78), .data_i_79_(subbytes_data_i_79), .data_i_80_(subbytes_data_i_80), .data_i_81_(subbytes_data_i_81), .data_i_82_(subbytes_data_i_82), .data_i_83_(subbytes_data_i_83), .data_i_84_(subbytes_data_i_84), .data_i_85_(subbytes_data_i_85), .data_i_86_(subbytes_data_i_86), .data_i_87_(subbytes_data_i_87), .data_i_88_(subbytes_data_i_88), .data_i_89_(subbytes_data_i_89), .data_i_90_(subbytes_data_i_90), .data_i_91_(subbytes_data_i_91), .data_i_92_(subbytes_data_i_92), .data_i_93_(subbytes_data_i_93), .data_i_94_(subbytes_data_i_94), .data_i_95_(subbytes_data_i_95), .data_i_96_(subbytes_data_i_96), .data_i_97_(subbytes_data_i_97), .data_i_98_(subbytes_data_i_98), .data_i_99_(subbytes_data_i_99), .data_i_100_(subbytes_data_i_100), .data_i_101_(subbytes_data_i_101), .data_i_102_(subbytes_data_i_102), .data_i_103_(subbytes_data_i_103), .data_i_104_(subbytes_data_i_104), .data_i_105_(subbytes_data_i_105), .data_i_106_(subbytes_data_i_106), .data_i_107_(subbytes_data_i_107), .data_i_108_(subbytes_data_i_108), .data_i_109_(subbytes_data_i_109), .data_i_110_(subbytes_data_i_110), .data_i_111_(subbytes_data_i_111), .data_i_112_(subbytes_data_i_112), .data_i_113_(subbytes_data_i_113), .data_i_114_(subbytes_data_i_114), .data_i_115_(subbytes_data_i_115), .data_i_116_(subbytes_data_i_116), .data_i_117_(subbytes_data_i_117), .data_i_118_(subbytes_data_i_118), .data_i_119_(subbytes_data_i_119), .data_i_120_(subbytes_data_i_120), .data_i_121_(subbytes_data_i_121), .data_i_122_(subbytes_data_i_122), .data_i_123_(subbytes_data_i_123), .data_i_124_(subbytes_data_i_124), .data_i_125_(subbytes_data_i_125), .data_i_126_(subbytes_data_i_126), .data_i_127_(subbytes_data_i_127), .data_o_0_(subbytes_data_o_0), .data_o_1_(subbytes_data_o_1), .data_o_2_(subbytes_data_o_2), .data_o_3_(subbytes_data_o_3), .data_o_4_(subbytes_data_o_4), .data_o_5_(subbytes_data_o_5), .data_o_6_(subbytes_data_o_6), .data_o_7_(subbytes_data_o_7), .data_o_8_(subbytes_data_o_8), .data_o_9_(subbytes_data_o_9), .data_o_10_(subbytes_data_o_10), .data_o_11_(subbytes_data_o_11), .data_o_12_(subbytes_data_o_12), .data_o_13_(subbytes_data_o_13), .data_o_14_(subbytes_data_o_14), .data_o_15_(subbytes_data_o_15), .data_o_16_(subbytes_data_o_16), .data_o_17_(subbytes_data_o_17), .data_o_18_(subbytes_data_o_18), .data_o_19_(subbytes_data_o_19), .data_o_20_(subbytes_data_o_20), .data_o_21_(subbytes_data_o_21), .data_o_22_(subbytes_data_o_22), .data_o_23_(subbytes_data_o_23), .data_o_24_(subbytes_data_o_24), .data_o_25_(subbytes_data_o_25), .data_o_26_(subbytes_data_o_26), .data_o_27_(subbytes_data_o_27), .data_o_28_(subbytes_data_o_28), .data_o_29_(subbytes_data_o_29), .data_o_30_(subbytes_data_o_30), .data_o_31_(subbytes_data_o_31), .data_o_32_(subbytes_data_o_32), .data_o_33_(subbytes_data_o_33), .data_o_34_(subbytes_data_o_34), .data_o_35_(subbytes_data_o_35), .data_o_36_(subbytes_data_o_36), .data_o_37_(subbytes_data_o_37), .data_o_38_(subbytes_data_o_38), .data_o_39_(subbytes_data_o_39), .data_o_40_(subbytes_data_o_40), .data_o_41_(subbytes_data_o_41), .data_o_42_(subbytes_data_o_42), .data_o_43_(subbytes_data_o_43), .data_o_44_(subbytes_data_o_44), .data_o_45_(subbytes_data_o_45), .data_o_46_(subbytes_data_o_46), .data_o_47_(subbytes_data_o_47), .data_o_48_(subbytes_data_o_48), .data_o_49_(subbytes_data_o_49), .data_o_50_(subbytes_data_o_50), .data_o_51_(subbytes_data_o_51), .data_o_52_(subbytes_data_o_52), .data_o_53_(subbytes_data_o_53), .data_o_54_(subbytes_data_o_54), .data_o_55_(subbytes_data_o_55), .data_o_56_(subbytes_data_o_56), .data_o_57_(subbytes_data_o_57), .data_o_58_(subbytes_data_o_58), .data_o_59_(subbytes_data_o_59), .data_o_60_(subbytes_data_o_60), .data_o_61_(subbytes_data_o_61), .data_o_62_(subbytes_data_o_62), .data_o_63_(subbytes_data_o_63), .data_o_64_(subbytes_data_o_64), .data_o_65_(subbytes_data_o_65), .data_o_66_(subbytes_data_o_66), .data_o_67_(subbytes_data_o_67), .data_o_68_(subbytes_data_o_68), .data_o_69_(subbytes_data_o_69), .data_o_70_(subbytes_data_o_70), .data_o_71_(subbytes_data_o_71), .data_o_72_(subbytes_data_o_72), .data_o_73_(subbytes_data_o_73), .data_o_74_(subbytes_data_o_74), .data_o_75_(subbytes_data_o_75), .data_o_76_(subbytes_data_o_76), .data_o_77_(subbytes_data_o_77), .data_o_78_(subbytes_data_o_78), .data_o_79_(subbytes_data_o_79), .data_o_80_(subbytes_data_o_80), .data_o_81_(subbytes_data_o_81), .data_o_82_(subbytes_data_o_82), .data_o_83_(subbytes_data_o_83), .data_o_84_(subbytes_data_o_84), .data_o_85_(subbytes_data_o_85), .data_o_86_(subbytes_data_o_86), .data_o_87_(subbytes_data_o_87), .data_o_88_(subbytes_data_o_88), .data_o_89_(subbytes_data_o_89), .data_o_90_(subbytes_data_o_90), .data_o_91_(subbytes_data_o_91), .data_o_92_(subbytes_data_o_92), .data_o_93_(subbytes_data_o_93), .data_o_94_(subbytes_data_o_94), .data_o_95_(subbytes_data_o_95), .data_o_96_(subbytes_data_o_96), .data_o_97_(subbytes_data_o_97), .data_o_98_(subbytes_data_o_98), .data_o_99_(subbytes_data_o_99), .data_o_100_(subbytes_data_o_100), .data_o_101_(subbytes_data_o_101), .data_o_102_(subbytes_data_o_102), .data_o_103_(subbytes_data_o_103), .data_o_104_(subbytes_data_o_104), .data_o_105_(subbytes_data_o_105), .data_o_106_(subbytes_data_o_106), .data_o_107_(subbytes_data_o_107), .data_o_108_(subbytes_data_o_108), .data_o_109_(subbytes_data_o_109), .data_o_110_(subbytes_data_o_110), .data_o_111_(subbytes_data_o_111), .data_o_112_(subbytes_data_o_112), .data_o_113_(subbytes_data_o_113), .data_o_114_(subbytes_data_o_114), .data_o_115_(subbytes_data_o_115), .data_o_116_(subbytes_data_o_116), .data_o_117_(subbytes_data_o_117), .data_o_118_(subbytes_data_o_118), .data_o_119_(subbytes_data_o_119), .data_o_120_(subbytes_data_o_120), .data_o_121_(subbytes_data_o_121), .data_o_122_(subbytes_data_o_122), .data_o_123_(subbytes_data_o_123), .data_o_124_(subbytes_data_o_124), .data_o_125_(subbytes_data_o_125), .data_o_126_(subbytes_data_o_126), .data_o_127_(subbytes_data_o_127), .decrypt_i(decrypt_i), .ready_o(subbytes_ready_o), .reset(reset), .sbox_data_i_0_(n4224), .sbox_data_i_1_(n4261), .sbox_data_i_2_(n4227), .sbox_data_i_3_(n4225), .sbox_data_i_4_(n4223), .sbox_data_i_5_(n4237), .sbox_data_i_6_(n4274), .sbox_data_i_7_(n4269), .sbox_data_o_0_(subbytes_sbox_data_o_0), .sbox_data_o_1_(subbytes_sbox_data_o_1), .sbox_data_o_2_(subbytes_sbox_data_o_2), .sbox_data_o_3_(subbytes_sbox_data_o_3), .sbox_data_o_4_(subbytes_sbox_data_o_4), .sbox_data_o_5_(subbytes_sbox_data_o_5), .sbox_data_o_6_(subbytes_sbox_data_o_6), .sbox_data_o_7_(subbytes_sbox_data_o_7), .sbox_decrypt_o(subbytes_sbox_decrypt_o), .start_i(subbytes_start_i));
endmodule

module subbytes (clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_i_8_, data_i_9_, data_i_10_, data_i_11_, data_i_12_, data_i_13_, data_i_14_, data_i_15_, data_i_16_, data_i_17_, data_i_18_, data_i_19_, data_i_20_, data_i_21_, data_i_22_, data_i_23_, data_i_24_, data_i_25_, data_i_26_, data_i_27_, data_i_28_, data_i_29_, data_i_30_, data_i_31_, data_i_32_, data_i_33_, data_i_34_, data_i_35_, data_i_36_, data_i_37_, data_i_38_, data_i_39_, data_i_40_, data_i_41_, data_i_42_, data_i_43_, data_i_44_, data_i_45_, data_i_46_, data_i_47_, data_i_48_, data_i_49_, data_i_50_, data_i_51_, data_i_52_, data_i_53_, data_i_54_, data_i_55_, data_i_56_, data_i_57_, data_i_58_, data_i_59_, data_i_60_, data_i_61_, data_i_62_, data_i_63_, data_i_64_, data_i_65_, data_i_66_, data_i_67_, data_i_68_, data_i_69_, data_i_70_, data_i_71_, data_i_72_, data_i_73_, data_i_74_, data_i_75_, data_i_76_, data_i_77_, data_i_78_, data_i_79_, data_i_80_, data_i_81_, data_i_82_, data_i_83_, data_i_84_, data_i_85_, data_i_86_, data_i_87_, data_i_88_, data_i_89_, data_i_90_, data_i_91_, data_i_92_, data_i_93_, data_i_94_, data_i_95_, data_i_96_, data_i_97_, data_i_98_, data_i_99_, data_i_100_, data_i_101_, data_i_102_, data_i_103_, data_i_104_, data_i_105_, data_i_106_, data_i_107_, data_i_108_, data_i_109_, data_i_110_, data_i_111_, data_i_112_, data_i_113_, data_i_114_, data_i_115_, data_i_116_, data_i_117_, data_i_118_, data_i_119_, data_i_120_, data_i_121_, data_i_122_, data_i_123_, data_i_124_, data_i_125_, data_i_126_, data_i_127_, data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_, data_o_32_, data_o_33_, data_o_34_, data_o_35_, data_o_36_, data_o_37_, data_o_38_, data_o_39_, data_o_40_, data_o_41_, data_o_42_, data_o_43_, data_o_44_, data_o_45_, data_o_46_, data_o_47_, data_o_48_, data_o_49_, data_o_50_, data_o_51_, data_o_52_, data_o_53_, data_o_54_, data_o_55_, data_o_56_, data_o_57_, data_o_58_, data_o_59_, data_o_60_, data_o_61_, data_o_62_, data_o_63_, data_o_64_, data_o_65_, data_o_66_, data_o_67_, data_o_68_, data_o_69_, data_o_70_, data_o_71_, data_o_72_, data_o_73_, data_o_74_, data_o_75_, data_o_76_, data_o_77_, data_o_78_, data_o_79_, data_o_80_, data_o_81_, data_o_82_, data_o_83_, data_o_84_, data_o_85_, data_o_86_, data_o_87_, data_o_88_, data_o_89_, data_o_90_, data_o_91_, data_o_92_, data_o_93_, data_o_94_, data_o_95_, data_o_96_, data_o_97_, data_o_98_, data_o_99_, data_o_100_, data_o_101_, data_o_102_, data_o_103_, data_o_104_, data_o_105_, data_o_106_, data_o_107_, data_o_108_, data_o_109_, data_o_110_, data_o_111_, data_o_112_, data_o_113_, data_o_114_, data_o_115_, data_o_116_, data_o_117_, data_o_118_, data_o_119_, data_o_120_, data_o_121_, data_o_122_, data_o_123_, data_o_124_, data_o_125_, data_o_126_, data_o_127_, decrypt_i, ready_o, reset, sbox_data_i_0_, sbox_data_i_1_, sbox_data_i_2_, sbox_data_i_3_, sbox_data_i_4_, sbox_data_i_5_, sbox_data_i_6_, sbox_data_i_7_, sbox_data_o_0_, sbox_data_o_1_, sbox_data_o_2_, sbox_data_o_3_, sbox_data_o_4_, sbox_data_o_5_, sbox_data_o_6_, sbox_data_o_7_, sbox_decrypt_o, start_i);
input clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_i_8_, data_i_9_, data_i_10_, data_i_11_, data_i_12_, data_i_13_, data_i_14_, data_i_15_, data_i_16_, data_i_17_, data_i_18_, data_i_19_, data_i_20_, data_i_21_, data_i_22_, data_i_23_, data_i_24_, data_i_25_, data_i_26_, data_i_27_, data_i_28_, data_i_29_, data_i_30_, data_i_31_, data_i_32_, data_i_33_, data_i_34_, data_i_35_, data_i_36_, data_i_37_, data_i_38_, data_i_39_, data_i_40_, data_i_41_, data_i_42_, data_i_43_, data_i_44_, data_i_45_, data_i_46_, data_i_47_, data_i_48_, data_i_49_, data_i_50_, data_i_51_, data_i_52_, data_i_53_, data_i_54_, data_i_55_, data_i_56_, data_i_57_, data_i_58_, data_i_59_, data_i_60_, data_i_61_, data_i_62_, data_i_63_, data_i_64_, data_i_65_, data_i_66_, data_i_67_, data_i_68_, data_i_69_, data_i_70_, data_i_71_, data_i_72_, data_i_73_, data_i_74_, data_i_75_, data_i_76_, data_i_77_, data_i_78_, data_i_79_, data_i_80_, data_i_81_, data_i_82_, data_i_83_, data_i_84_, data_i_85_, data_i_86_, data_i_87_, data_i_88_, data_i_89_, data_i_90_, data_i_91_, data_i_92_, data_i_93_, data_i_94_, data_i_95_, data_i_96_, data_i_97_, data_i_98_, data_i_99_, data_i_100_, data_i_101_, data_i_102_, data_i_103_, data_i_104_, data_i_105_, data_i_106_, data_i_107_, data_i_108_, data_i_109_, data_i_110_, data_i_111_, data_i_112_, data_i_113_, data_i_114_, data_i_115_, data_i_116_, data_i_117_, data_i_118_, data_i_119_, data_i_120_, data_i_121_, data_i_122_, data_i_123_, data_i_124_, data_i_125_, data_i_126_, data_i_127_, decrypt_i, reset, sbox_data_i_0_, sbox_data_i_1_, sbox_data_i_2_, sbox_data_i_3_, sbox_data_i_4_, sbox_data_i_5_, sbox_data_i_6_, sbox_data_i_7_, start_i;
output data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_, data_o_32_, data_o_33_, data_o_34_, data_o_35_, data_o_36_, data_o_37_, data_o_38_, data_o_39_, data_o_40_, data_o_41_, data_o_42_, data_o_43_, data_o_44_, data_o_45_, data_o_46_, data_o_47_, data_o_48_, data_o_49_, data_o_50_, data_o_51_, data_o_52_, data_o_53_, data_o_54_, data_o_55_, data_o_56_, data_o_57_, data_o_58_, data_o_59_, data_o_60_, data_o_61_, data_o_62_, data_o_63_, data_o_64_, data_o_65_, data_o_66_, data_o_67_, data_o_68_, data_o_69_, data_o_70_, data_o_71_, data_o_72_, data_o_73_, data_o_74_, data_o_75_, data_o_76_, data_o_77_, data_o_78_, data_o_79_, data_o_80_, data_o_81_, data_o_82_, data_o_83_, data_o_84_, data_o_85_, data_o_86_, data_o_87_, data_o_88_, data_o_89_, data_o_90_, data_o_91_, data_o_92_, data_o_93_, data_o_94_, data_o_95_, data_o_96_, data_o_97_, data_o_98_, data_o_99_, data_o_100_, data_o_101_, data_o_102_, data_o_103_, data_o_104_, data_o_105_, data_o_106_, data_o_107_, data_o_108_, data_o_109_, data_o_110_, data_o_111_, data_o_112_, data_o_113_, data_o_114_, data_o_115_, data_o_116_, data_o_117_, data_o_118_, data_o_119_, data_o_120_, data_o_121_, data_o_122_, data_o_123_, data_o_124_, data_o_125_, data_o_126_, data_o_127_, ready_o, sbox_data_o_0_, sbox_data_o_1_, sbox_data_o_2_, sbox_data_o_3_, sbox_data_o_4_, sbox_data_o_5_, sbox_data_o_6_, sbox_data_o_7_, sbox_decrypt_o;

sg13g2_nand3_1 U1 (.A(n317), .B(n727), .C(n726), .Y(n741));
sg13g2_nand3_1 U2 (.A(n321), .B(n648), .C(n647), .Y(n668));
sg13g2_inv_4 U3 (.A(n790), .Y(n584));
sg13g2_nand2_2 U4 (.A(data_i_127_), .B(n4), .Y(n3));
sg13g2_o21ai_1 U5 (.A1(n46), .A2(n45), .B1(n47), .Y(n477));
sg13g2_o21ai_1 U6 (.A1(n51), .A2(n45), .B1(n260), .Y(n525));
sg13g2_nand2_2 U7 (.A(data_i_126_), .B(n4), .Y(n6));
sg13g2_nand2_2 U8 (.A(N32), .B(N31), .Y(n598));
sg13g2_o21ai_1 U9 (.A1(n197), .A2(n45), .B1(n405), .Y(n459));
sg13g2_nand2_2 U10 (.A(data_i_125_), .B(n4), .Y(n8));
sg13g2_nor2_2 U11 (.A(n590), .B(N31), .Y(n600));
sg13g2_o21ai_1 U12 (.A1(n9), .A2(n1), .B1(n10), .Y(sbox_data_o_4_));
sg13g2_nand2_2 U13 (.A(data_i_124_), .B(n4), .Y(n10));
sg13g2_inv_4 U14 (.A(N127), .Y(n9));
sg13g2_o21ai_1 U15 (.A1(n194), .A2(n45), .B1(n195), .Y(n507));
sg13g2_nor2_2 U16 (.A(N31), .B(N32), .Y(n596));
sg13g2_o21ai_1 U17 (.A1(n7), .A2(n1), .B1(n8), .Y(sbox_data_o_5_));
sg13g2_inv_4 U18 (.A(N126), .Y(n7));
sg13g2_nand2_2 U19 (.A(data_i_122_), .B(n4), .Y(n14));
sg13g2_inv_4 U20 (.A(N129), .Y(n13));
sg13g2_o21ai_1 U21 (.A1(n189), .A2(n45), .B1(n401), .Y(n457));
sg13g2_nand2_2 U22 (.A(data_i_121_), .B(n4), .Y(n16));
sg13g2_o21ai_1 U23 (.A1(n693), .A2(n692), .B1(n691), .Y(N128));
sg13g2_o21ai_1 U24 (.A1(n17), .A2(n1), .B1(n18), .Y(sbox_data_o_0_));
sg13g2_nand2_2 U25 (.A(data_i_120_), .B(n4), .Y(n18));
sg13g2_o21ai_1 U26 (.A1(n186), .A2(n45), .B1(n187), .Y(n505));
sg13g2_o21ai_1 U27 (.A1(n13), .A2(n1), .B1(n14), .Y(sbox_data_o_2_));
sg13g2_nand3_1 U28 (.A(n588), .B(n751), .C(n750), .Y(n766));
sg13g2_a21oi_2 U29 (.A1(sbox_data_i_3_), .A2(n25), .B1(n26), .Y(n24));
sg13g2_nor2_2 U30 (.A(n27), .B(n28), .Y(n26));
sg13g2_nand2_2 U31 (.A(data_o_51_), .B(n29), .Y(n23));
sg13g2_nand3_1 U32 (.A(n747), .B(n746), .C(n745), .Y(n767));
sg13g2_a21oi_2 U33 (.A1(sbox_data_i_2_), .A2(n25), .B1(n33), .Y(n32));
sg13g2_nor2_2 U34 (.A(n27), .B(n34), .Y(n33));
sg13g2_nand2_2 U35 (.A(data_o_50_), .B(n29), .Y(n31));
sg13g2_nand3_1 U36 (.A(n807), .B(n673), .C(n672), .Y(n693));
sg13g2_a21oi_2 U37 (.A1(sbox_data_i_1_), .A2(n25), .B1(n38), .Y(n37));
sg13g2_nor2_2 U38 (.A(n27), .B(n39), .Y(n38));
sg13g2_nand2_2 U39 (.A(data_o_49_), .B(n29), .Y(n36));
sg13g2_nand3_1 U40 (.A(n808), .B(n678), .C(n677), .Y(n692));
sg13g2_a21oi_2 U41 (.A1(sbox_data_i_0_), .A2(n25), .B1(n43), .Y(n42));
sg13g2_nor2_2 U42 (.A(n27), .B(n44), .Y(n43));
sg13g2_nand2_2 U43 (.A(data_o_48_), .B(n29), .Y(n41));
sg13g2_o21ai_1 U44 (.A1(n181), .A2(n45), .B1(n397), .Y(n455));
sg13g2_a21oi_2 U45 (.A1(sbox_data_i_7_), .A2(n48), .B1(n49), .Y(n47));
sg13g2_nor2_2 U46 (.A(n50), .B(n51), .Y(n49));
sg13g2_o21ai_1 U47 (.A1(n587), .A2(n52), .B1(n53), .Y(n478));
sg13g2_a21oi_2 U48 (.A1(sbox_data_i_6_), .A2(n48), .B1(n54), .Y(n53));
sg13g2_nor2_2 U49 (.A(n50), .B(n55), .Y(n54));
sg13g2_o21ai_1 U50 (.A1(n45), .A2(n56), .B1(n57), .Y(n479));
sg13g2_a21oi_2 U51 (.A1(sbox_data_i_5_), .A2(n48), .B1(n58), .Y(n57));
sg13g2_nor2_2 U52 (.A(n50), .B(n59), .Y(n58));
sg13g2_o21ai_1 U53 (.A1(n587), .A2(n60), .B1(n61), .Y(n480));
sg13g2_a21oi_2 U54 (.A1(sbox_data_i_4_), .A2(n48), .B1(n62), .Y(n61));
sg13g2_nor2_2 U55 (.A(n50), .B(n63), .Y(n62));
sg13g2_o21ai_1 U56 (.A1(n45), .A2(n64), .B1(n65), .Y(n481));
sg13g2_a21oi_2 U57 (.A1(n48), .A2(sbox_data_i_3_), .B1(n66), .Y(n65));
sg13g2_nor2_2 U58 (.A(n50), .B(n67), .Y(n66));
sg13g2_o21ai_1 U59 (.A1(n587), .A2(n68), .B1(n69), .Y(n482));
sg13g2_a21oi_2 U60 (.A1(n48), .A2(sbox_data_i_2_), .B1(n70), .Y(n69));
sg13g2_nor2_2 U61 (.A(n50), .B(n71), .Y(n70));
sg13g2_o21ai_1 U62 (.A1(n45), .A2(n72), .B1(n73), .Y(n483));
sg13g2_a21oi_2 U63 (.A1(n48), .A2(sbox_data_i_1_), .B1(n74), .Y(n73));
sg13g2_nor2_2 U64 (.A(n50), .B(n75), .Y(n74));
sg13g2_o21ai_1 U65 (.A1(n587), .A2(n76), .B1(n77), .Y(n484));
sg13g2_a21oi_2 U66 (.A1(n48), .A2(sbox_data_i_0_), .B1(n78), .Y(n77));
sg13g2_nor2_2 U67 (.A(n50), .B(n79), .Y(n78));
sg13g2_nand2_2 U68 (.A(n80), .B(n587), .Y(n50));
sg13g2_inv_4 U69 (.A(n80), .Y(n48));
sg13g2_nand2_2 U70 (.A(n81), .B(n82), .Y(n80));
sg13g2_nand3_1 U71 (.A(n809), .B(n603), .C(n602), .Y(n617));
sg13g2_a21oi_2 U72 (.A1(n86), .A2(sbox_data_i_7_), .B1(n87), .Y(n85));
sg13g2_nor2_2 U73 (.A(n88), .B(n89), .Y(n87));
sg13g2_nand2_2 U74 (.A(data_o_103_), .B(n29), .Y(n84));
sg13g2_nand3_1 U75 (.A(n810), .B(n594), .C(n593), .Y(n618));
sg13g2_a21oi_2 U76 (.A1(n86), .A2(sbox_data_i_6_), .B1(n93), .Y(n92));
sg13g2_nor2_2 U77 (.A(n88), .B(n94), .Y(n93));
sg13g2_nand2_2 U78 (.A(data_o_102_), .B(n29), .Y(n91));
sg13g2_nand3_1 U79 (.A(n697), .B(n811), .C(n322), .Y(n717));
sg13g2_a21oi_2 U80 (.A1(n86), .A2(sbox_data_i_5_), .B1(n98), .Y(n97));
sg13g2_nor2_2 U81 (.A(n88), .B(n99), .Y(n98));
sg13g2_nand2_2 U82 (.A(data_o_101_), .B(n29), .Y(n96));
sg13g2_nand3_1 U83 (.A(n812), .B(n702), .C(n701), .Y(n716));
sg13g2_a21oi_2 U84 (.A1(n86), .A2(sbox_data_i_4_), .B1(n103), .Y(n102));
sg13g2_nor2_2 U85 (.A(n88), .B(n104), .Y(n103));
sg13g2_nand2_2 U86 (.A(data_o_100_), .B(n29), .Y(n101));
sg13g2_nand3_1 U87 (.A(n772), .B(n813), .C(n773), .Y(n802));
sg13g2_a21oi_2 U88 (.A1(n86), .A2(sbox_data_i_3_), .B1(n108), .Y(n107));
sg13g2_nor2_2 U89 (.A(n88), .B(n109), .Y(n108));
sg13g2_nand2_2 U90 (.A(data_o_99_), .B(n29), .Y(n106));
sg13g2_a21oi_1 U91 (.A1(n814), .A2(n794), .B1(n793), .Y(n796));
sg13g2_o21ai_1 U92 (.A1(n767), .A2(n766), .B1(n765), .Y(N125));
sg13g2_nor2_2 U93 (.A(n88), .B(n114), .Y(n113));
sg13g2_nand2_2 U94 (.A(data_o_98_), .B(n29), .Y(n111));
sg13g2_nand3_1 U95 (.A(N33), .B(n815), .C(n777), .Y(n801));
sg13g2_a21oi_2 U96 (.A1(n86), .A2(sbox_data_i_1_), .B1(n118), .Y(n117));
sg13g2_nor2_2 U97 (.A(n88), .B(n119), .Y(n118));
sg13g2_nand2_2 U98 (.A(data_o_97_), .B(n29), .Y(n116));
sg13g2_nand3_1 U99 (.A(n816), .B(n623), .C(n622), .Y(n643));
sg13g2_a21oi_2 U100 (.A1(n86), .A2(sbox_data_i_0_), .B1(n123), .Y(n122));
sg13g2_nor2_2 U101 (.A(n88), .B(n124), .Y(n123));
sg13g2_nand2_2 U102 (.A(n125), .B(n587), .Y(n88));
sg13g2_inv_4 U103 (.A(n125), .Y(n86));
sg13g2_nand2_2 U104 (.A(n126), .B(n127), .Y(n125));
sg13g2_nand2_2 U105 (.A(data_o_96_), .B(n29), .Y(n121));
sg13g2_nand3_1 U106 (.A(n817), .B(n628), .C(n627), .Y(n642));
sg13g2_a21oi_2 U107 (.A1(n131), .A2(sbox_data_i_7_), .B1(n132), .Y(n130));
sg13g2_nor2_2 U108 (.A(n133), .B(n134), .Y(n132));
sg13g2_nand2_2 U109 (.A(data_o_23_), .B(n29), .Y(n129));
sg13g2_nand3_1 U110 (.A(n818), .B(n722), .C(n721), .Y(n742));
sg13g2_a21oi_2 U111 (.A1(n131), .A2(sbox_data_i_6_), .B1(n138), .Y(n137));
sg13g2_nor2_2 U112 (.A(n133), .B(n139), .Y(n138));
sg13g2_nand2_2 U113 (.A(data_o_22_), .B(n29), .Y(n136));
sg13g2_nand3_1 U114 (.A(n819), .B(n653), .C(n652), .Y(n667));
sg13g2_a21oi_2 U115 (.A1(n131), .A2(sbox_data_i_5_), .B1(n143), .Y(n142));
sg13g2_nor2_2 U116 (.A(n133), .B(n144), .Y(n143));
sg13g2_nand2_2 U117 (.A(data_o_21_), .B(n29), .Y(n141));
sg13g2_nand3_1 U118 (.A(n440), .B(n820), .C(n439), .Y(n472));
sg13g2_a21oi_2 U119 (.A1(n131), .A2(sbox_data_i_4_), .B1(n148), .Y(n147));
sg13g2_nor2_2 U120 (.A(n133), .B(n149), .Y(n148));
sg13g2_nand2_2 U121 (.A(data_o_20_), .B(n29), .Y(n146));
sg13g2_nand3_1 U122 (.A(n437), .B(n821), .C(n436), .Y(n471));
sg13g2_a21oi_2 U123 (.A1(n131), .A2(sbox_data_i_3_), .B1(n152), .Y(n151));
sg13g2_nor2_2 U124 (.A(n153), .B(n133), .Y(n152));
sg13g2_nand2_2 U125 (.A(data_o_19_), .B(n29), .Y(n150));
sg13g2_nand3_1 U126 (.A(n434), .B(n822), .C(n433), .Y(n470));
sg13g2_nand3_1 U127 (.A(n431), .B(n823), .C(n430), .Y(n469));
sg13g2_a21oi_2 U128 (.A1(n131), .A2(sbox_data_i_2_), .B1(n156), .Y(n155));
sg13g2_nor2_2 U129 (.A(n157), .B(n133), .Y(n156));
sg13g2_nand2_2 U130 (.A(data_o_18_), .B(n29), .Y(n154));
sg13g2_nand3_1 U131 (.A(n388), .B(n824), .C(n387), .Y(n452));
sg13g2_nand3_1 U132 (.A(n385), .B(n825), .C(n384), .Y(n451));
sg13g2_a21oi_2 U133 (.A1(n131), .A2(sbox_data_i_1_), .B1(n160), .Y(n159));
sg13g2_nor2_2 U134 (.A(n161), .B(n133), .Y(n160));
sg13g2_nand2_2 U135 (.A(data_o_17_), .B(n29), .Y(n158));
sg13g2_nand3_1 U136 (.A(n382), .B(n826), .C(n381), .Y(n450));
sg13g2_nand3_1 U137 (.A(n379), .B(n827), .C(n378), .Y(n449));
sg13g2_a21oi_2 U138 (.A1(n131), .A2(sbox_data_i_0_), .B1(n164), .Y(n163));
sg13g2_nor2_2 U139 (.A(n165), .B(n133), .Y(n164));
sg13g2_nand2_2 U140 (.A(n166), .B(n587), .Y(n133));
sg13g2_inv_4 U141 (.A(n166), .Y(n131));
sg13g2_nand2_2 U142 (.A(n126), .B(n167), .Y(n166));
sg13g2_nand2_2 U143 (.A(data_o_16_), .B(n29), .Y(n162));
sg13g2_nand3_1 U144 (.A(n375), .B(n828), .C(n374), .Y(n448));
sg13g2_mux2_2 U145 (.A0(sbox_data_i_7_), .A1(data_o_31_), .S(n304), .X(n547));
sg13g2_a21oi_2 U146 (.A1(n170), .A2(sbox_data_i_7_), .B1(n171), .Y(n169));
sg13g2_nor2_2 U147 (.A(n172), .B(n173), .Y(n171));
sg13g2_o21ai_1 U148 (.A1(n587), .A2(n174), .B1(n175), .Y(n502));
sg13g2_a21oi_2 U149 (.A1(n170), .A2(sbox_data_i_6_), .B1(n176), .Y(n175));
sg13g2_nor2_2 U150 (.A(n172), .B(n177), .Y(n176));
sg13g2_nand3_1 U151 (.A(n371), .B(n829), .C(n370), .Y(n447));
sg13g2_a21oi_2 U152 (.A1(n170), .A2(sbox_data_i_5_), .B1(n180), .Y(n179));
sg13g2_nor2_2 U153 (.A(n172), .B(n181), .Y(n180));
sg13g2_o21ai_1 U154 (.A1(n587), .A2(n182), .B1(n183), .Y(n504));
sg13g2_a21oi_2 U155 (.A1(n170), .A2(sbox_data_i_4_), .B1(n184), .Y(n183));
sg13g2_nor2_2 U156 (.A(n172), .B(n185), .Y(n184));
sg13g2_o21ai_1 U157 (.A1(n119), .A2(n203), .B1(n218), .Y(n515));
sg13g2_a21oi_2 U158 (.A1(n170), .A2(sbox_data_i_3_), .B1(n188), .Y(n187));
sg13g2_nor2_2 U159 (.A(n172), .B(n189), .Y(n188));
sg13g2_o21ai_1 U160 (.A1(n587), .A2(n190), .B1(n191), .Y(n506));
sg13g2_a21oi_2 U161 (.A1(n170), .A2(sbox_data_i_2_), .B1(n192), .Y(n191));
sg13g2_nor2_2 U162 (.A(n172), .B(n193), .Y(n192));
sg13g2_o21ai_1 U163 (.A1(n178), .A2(n45), .B1(n179), .Y(n503));
sg13g2_a21oi_2 U164 (.A1(n170), .A2(sbox_data_i_1_), .B1(n196), .Y(n195));
sg13g2_nor2_2 U165 (.A(n172), .B(n197), .Y(n196));
sg13g2_o21ai_1 U166 (.A1(n587), .A2(n198), .B1(n199), .Y(n508));
sg13g2_a21oi_2 U167 (.A1(n170), .A2(sbox_data_i_0_), .B1(n200), .Y(n199));
sg13g2_nor2_2 U168 (.A(n172), .B(n201), .Y(n200));
sg13g2_nand2_2 U169 (.A(n202), .B(n587), .Y(n172));
sg13g2_inv_4 U170 (.A(n202), .Y(n170));
sg13g2_nand2_2 U171 (.A(n126), .B(n81), .Y(n202));
sg13g2_o21ai_1 U172 (.A1(n203), .A2(n89), .B1(n204), .Y(n509));
sg13g2_a21oi_2 U173 (.A1(sbox_data_i_7_), .A2(n205), .B1(n206), .Y(n204));
sg13g2_nor2_2 U174 (.A(n83), .B(n207), .Y(n206));
sg13g2_nand3_1 U175 (.A(n367), .B(n830), .C(n366), .Y(n446));
sg13g2_o21ai_1 U176 (.A1(n203), .A2(n94), .B1(n208), .Y(n510));
sg13g2_a21oi_2 U177 (.A1(sbox_data_i_6_), .A2(n205), .B1(n209), .Y(n208));
sg13g2_nor2_2 U178 (.A(n90), .B(n207), .Y(n209));
sg13g2_nand3_1 U179 (.A(n361), .B(n831), .C(n360), .Y(n445));
sg13g2_nand2_2 U180 (.A(n590), .B(N31), .Y(n595));
sg13g2_a21oi_2 U181 (.A1(sbox_data_i_5_), .A2(n205), .B1(n211), .Y(n210));
sg13g2_nor2_2 U182 (.A(n95), .B(n207), .Y(n211));
sg13g2_nand3_1 U183 (.A(n302), .B(n832), .C(n301), .Y(n540));
sg13g2_o21ai_1 U184 (.A1(n104), .A2(n203), .B1(n212), .Y(n512));
sg13g2_a21oi_2 U185 (.A1(sbox_data_i_4_), .A2(n205), .B1(n213), .Y(n212));
sg13g2_nor2_2 U186 (.A(n100), .B(n207), .Y(n213));
sg13g2_nand3_1 U187 (.A(n299), .B(n833), .C(n298), .Y(n539));
sg13g2_o21ai_1 U188 (.A1(n203), .A2(n109), .B1(n214), .Y(n513));
sg13g2_a21oi_2 U189 (.A1(sbox_data_i_3_), .A2(n205), .B1(n215), .Y(n214));
sg13g2_nor2_2 U190 (.A(n105), .B(n207), .Y(n215));
sg13g2_nand3_1 U191 (.A(n296), .B(n834), .C(n295), .Y(n538));
sg13g2_o21ai_1 U192 (.A1(n203), .A2(n114), .B1(n216), .Y(n514));
sg13g2_a21oi_2 U193 (.A1(sbox_data_i_2_), .A2(n205), .B1(n217), .Y(n216));
sg13g2_nor2_2 U194 (.A(n110), .B(n207), .Y(n217));
sg13g2_nand3_1 U195 (.A(n293), .B(n835), .C(n292), .Y(n537));
sg13g2_o21ai_1 U196 (.A1(n173), .A2(n45), .B1(n391), .Y(n453));
sg13g2_a21oi_2 U197 (.A1(sbox_data_i_1_), .A2(n205), .B1(n219), .Y(n218));
sg13g2_nor2_2 U198 (.A(n115), .B(n207), .Y(n219));
sg13g2_nand3_1 U199 (.A(n290), .B(n836), .C(n289), .Y(n536));
sg13g2_o21ai_1 U200 (.A1(n203), .A2(n124), .B1(n220), .Y(n516));
sg13g2_a21oi_2 U201 (.A1(sbox_data_i_0_), .A2(n205), .B1(n221), .Y(n220));
sg13g2_nor2_2 U202 (.A(n120), .B(n207), .Y(n221));
sg13g2_nand2_2 U203 (.A(n222), .B(n587), .Y(n207));
sg13g2_nand3_1 U204 (.A(n287), .B(n837), .C(n286), .Y(n535));
sg13g2_o21ai_1 U205 (.A1(n587), .A2(n223), .B1(n222), .Y(n205));
sg13g2_nand2_2 U206 (.A(n224), .B(n127), .Y(n222));
sg13g2_nand3_1 U207 (.A(n284), .B(n838), .C(n283), .Y(n534));
sg13g2_a21oi_2 U208 (.A1(n227), .A2(sbox_data_i_7_), .B1(n228), .Y(n226));
sg13g2_nor2_2 U209 (.A(n229), .B(n230), .Y(n228));
sg13g2_nand2_2 U210 (.A(data_o_119_), .B(n29), .Y(n225));
sg13g2_nand3_1 U211 (.A(n281), .B(n839), .C(n280), .Y(n533));
sg13g2_nand3_1 U212 (.A(n256), .B(n840), .C(n255), .Y(n524));
sg13g2_a21oi_2 U213 (.A1(n227), .A2(sbox_data_i_6_), .B1(n233), .Y(n232));
sg13g2_nor2_2 U214 (.A(n234), .B(n230), .Y(n233));
sg13g2_nand2_2 U215 (.A(data_o_118_), .B(n29), .Y(n231));
sg13g2_nand3_1 U216 (.A(n252), .B(n841), .C(n251), .Y(n523));
sg13g2_nand3_1 U217 (.A(n248), .B(n842), .C(n247), .Y(n522));
sg13g2_a21oi_2 U218 (.A1(n227), .A2(sbox_data_i_5_), .B1(n237), .Y(n236));
sg13g2_nor2_2 U219 (.A(n238), .B(n230), .Y(n237));
sg13g2_nand2_2 U220 (.A(data_o_117_), .B(n29), .Y(n235));
sg13g2_nand3_1 U221 (.A(n244), .B(n843), .C(n243), .Y(n521));
sg13g2_nand3_1 U222 (.A(n240), .B(n844), .C(n239), .Y(n520));
sg13g2_a21oi_2 U223 (.A1(n227), .A2(sbox_data_i_4_), .B1(n241), .Y(n240));
sg13g2_nor2_2 U224 (.A(n242), .B(n230), .Y(n241));
sg13g2_nand2_2 U225 (.A(data_o_116_), .B(n29), .Y(n239));
sg13g2_nand3_1 U226 (.A(n236), .B(n845), .C(n235), .Y(n519));
sg13g2_nand3_1 U227 (.A(n232), .B(n846), .C(n231), .Y(n518));
sg13g2_a21oi_2 U228 (.A1(n227), .A2(sbox_data_i_3_), .B1(n245), .Y(n244));
sg13g2_nor2_2 U229 (.A(n246), .B(n230), .Y(n245));
sg13g2_nand2_2 U230 (.A(data_o_115_), .B(n29), .Y(n243));
sg13g2_nand3_1 U231 (.A(n226), .B(n847), .C(n225), .Y(n517));
sg13g2_nand3_1 U232 (.A(n163), .B(n848), .C(n162), .Y(n500));
sg13g2_a21oi_2 U233 (.A1(n227), .A2(sbox_data_i_2_), .B1(n249), .Y(n248));
sg13g2_nor2_2 U234 (.A(n250), .B(n230), .Y(n249));
sg13g2_nand2_2 U235 (.A(data_o_114_), .B(n29), .Y(n247));
sg13g2_nand3_1 U236 (.A(n159), .B(n849), .C(n158), .Y(n499));
sg13g2_nand3_1 U237 (.A(n155), .B(n850), .C(n154), .Y(n498));
sg13g2_a21oi_2 U238 (.A1(n227), .A2(sbox_data_i_1_), .B1(n253), .Y(n252));
sg13g2_nor2_2 U239 (.A(n254), .B(n230), .Y(n253));
sg13g2_nand2_2 U240 (.A(data_o_113_), .B(n29), .Y(n251));
sg13g2_nand3_1 U241 (.A(n151), .B(n851), .C(n150), .Y(n497));
sg13g2_nand3_1 U242 (.A(n147), .B(n852), .C(n146), .Y(n496));
sg13g2_a21oi_2 U243 (.A1(n227), .A2(sbox_data_i_0_), .B1(n257), .Y(n256));
sg13g2_nor2_2 U244 (.A(n258), .B(n230), .Y(n257));
sg13g2_nand2_2 U245 (.A(n259), .B(n587), .Y(n230));
sg13g2_inv_4 U246 (.A(n259), .Y(n227));
sg13g2_nand2_2 U247 (.A(n224), .B(n167), .Y(n259));
sg13g2_nand2_2 U248 (.A(data_o_112_), .B(n29), .Y(n255));
sg13g2_nand3_1 U249 (.A(n142), .B(n853), .C(n141), .Y(n495));
sg13g2_o21ai_1 U250 (.A1(n15), .A2(n1), .B1(n16), .Y(sbox_data_o_1_));
sg13g2_a21oi_2 U251 (.A1(n261), .A2(sbox_data_i_7_), .B1(n262), .Y(n260));
sg13g2_nor2_2 U252 (.A(n46), .B(n263), .Y(n262));
sg13g2_nand3_1 U253 (.A(n137), .B(n854), .C(n136), .Y(n494));
sg13g2_nand3_1 U254 (.A(n130), .B(n855), .C(n129), .Y(n493));
sg13g2_o21ai_1 U255 (.A1(n587), .A2(n55), .B1(n264), .Y(n526));
sg13g2_a21oi_2 U256 (.A1(n261), .A2(sbox_data_i_6_), .B1(n265), .Y(n264));
sg13g2_nor2_2 U257 (.A(n52), .B(n263), .Y(n265));
sg13g2_nand3_1 U258 (.A(n122), .B(n856), .C(n121), .Y(n492));
sg13g2_nand3_1 U259 (.A(n117), .B(n857), .C(n116), .Y(n491));
sg13g2_o21ai_1 U260 (.A1(n45), .A2(n59), .B1(n266), .Y(n527));
sg13g2_a21oi_2 U261 (.A1(n261), .A2(sbox_data_i_5_), .B1(n267), .Y(n266));
sg13g2_nor2_2 U262 (.A(n56), .B(n263), .Y(n267));
sg13g2_nand3_1 U263 (.A(n112), .B(n858), .C(n111), .Y(n490));
sg13g2_nand3_1 U264 (.A(n107), .B(n859), .C(n106), .Y(n489));
sg13g2_o21ai_1 U265 (.A1(n587), .A2(n63), .B1(n268), .Y(n528));
sg13g2_a21oi_2 U266 (.A1(n261), .A2(sbox_data_i_4_), .B1(n269), .Y(n268));
sg13g2_nor2_2 U267 (.A(n60), .B(n263), .Y(n269));
sg13g2_nand3_1 U268 (.A(n102), .B(n860), .C(n101), .Y(n488));
sg13g2_nand3_1 U269 (.A(n97), .B(n861), .C(n96), .Y(n487));
sg13g2_o21ai_1 U270 (.A1(n45), .A2(n67), .B1(n270), .Y(n529));
sg13g2_a21oi_2 U271 (.A1(n261), .A2(sbox_data_i_3_), .B1(n271), .Y(n270));
sg13g2_nor2_2 U272 (.A(n64), .B(n263), .Y(n271));
sg13g2_nand3_1 U273 (.A(n92), .B(n862), .C(n91), .Y(n486));
sg13g2_nand3_1 U274 (.A(n85), .B(n863), .C(n84), .Y(n485));
sg13g2_o21ai_1 U275 (.A1(n587), .A2(n71), .B1(n272), .Y(n530));
sg13g2_a21oi_2 U276 (.A1(n261), .A2(sbox_data_i_2_), .B1(n273), .Y(n272));
sg13g2_nor2_2 U277 (.A(n68), .B(n263), .Y(n273));
sg13g2_nand3_1 U278 (.A(n42), .B(n864), .C(n41), .Y(n476));
sg13g2_nand3_1 U279 (.A(n37), .B(n865), .C(n36), .Y(n475));
sg13g2_o21ai_1 U280 (.A1(n45), .A2(n75), .B1(n274), .Y(n531));
sg13g2_a21oi_2 U281 (.A1(n261), .A2(sbox_data_i_1_), .B1(n275), .Y(n274));
sg13g2_nor2_2 U282 (.A(n72), .B(n263), .Y(n275));
sg13g2_nand3_1 U283 (.A(n32), .B(n866), .C(n31), .Y(n474));
sg13g2_nand3_1 U284 (.A(n24), .B(n867), .C(n23), .Y(n473));
sg13g2_o21ai_1 U285 (.A1(n587), .A2(n79), .B1(n276), .Y(n532));
sg13g2_a21oi_2 U286 (.A1(n261), .A2(sbox_data_i_0_), .B1(n277), .Y(n276));
sg13g2_nor2_2 U287 (.A(n76), .B(n263), .Y(n277));
sg13g2_nand2_2 U288 (.A(n278), .B(n587), .Y(n263));
sg13g2_nor2_1 U289 (.A(n595), .B(N30), .Y(n814));
sg13g2_inv_4 U290 (.A(n278), .Y(n261));
sg13g2_nand2_2 U291 (.A(n224), .B(n81), .Y(n278));
sg13g2_inv_1 U292 (.A(n21), .Y(n868));
sg13g2_or2_1 U293 (.A(data_i_31_), .B(n787), .X(n813));
sg13g2_nand2_2 U294 (.A(data_o_7_), .B(n45), .Y(n281));
sg13g2_nand2_2 U295 (.A(data_o_39_), .B(n29), .Y(n280));
sg13g2_nand2b_1 U296 (.A_N(data_i_7_), .B(n782), .Y(n815));
sg13g2_nand2_2 U297 (.A(data_o_6_), .B(n587), .Y(n284));
sg13g2_nand2_2 U298 (.A(data_o_38_), .B(n29), .Y(n283));
sg13g2_nand2b_1 U299 (.A_N(data_i_110_), .B(n795), .Y(n747));
sg13g2_nand2_2 U300 (.A(data_o_5_), .B(n45), .Y(n287));
sg13g2_nand2_2 U301 (.A(data_o_37_), .B(n29), .Y(n286));
sg13g2_or2_1 U302 (.A(n752), .B(data_i_102_), .X(n588));
sg13g2_nand2_2 U303 (.A(data_o_4_), .B(n587), .Y(n290));
sg13g2_nand2_2 U304 (.A(data_o_36_), .B(n29), .Y(n289));
sg13g2_nand2b_1 U305 (.A_N(data_i_109_), .B(n795), .Y(n818));
sg13g2_nand2_2 U306 (.A(data_o_3_), .B(n45), .Y(n293));
sg13g2_nand2_2 U307 (.A(data_o_35_), .B(n29), .Y(n292));
sg13g2_or2_1 U308 (.A(n752), .B(data_i_101_), .X(n317));
sg13g2_nand2_2 U309 (.A(data_o_2_), .B(n587), .Y(n296));
sg13g2_nand2_2 U310 (.A(data_o_34_), .B(n29), .Y(n295));
sg13g2_nand2b_1 U311 (.A_N(data_i_108_), .B(n795), .Y(n811));
sg13g2_nand2_2 U312 (.A(data_o_1_), .B(n587), .Y(n299));
sg13g2_nand2_2 U313 (.A(data_o_33_), .B(n29), .Y(n298));
sg13g2_or2_1 U314 (.A(n752), .B(data_i_100_), .X(n812));
sg13g2_nand2_2 U315 (.A(data_o_0_), .B(n587), .Y(n302));
sg13g2_nand2_2 U316 (.A(data_o_32_), .B(n29), .Y(n301));
sg13g2_o21ai_1 U317 (.A1(n303), .A2(n304), .B1(n305), .Y(n541));
sg13g2_nand2_2 U318 (.A(data_o_25_), .B(n304), .Y(n305));
sg13g2_o21ai_1 U319 (.A1(n306), .A2(n304), .B1(n307), .Y(n542));
sg13g2_nand2_2 U320 (.A(data_o_26_), .B(n304), .Y(n307));
sg13g2_o21ai_1 U321 (.A1(n308), .A2(n304), .B1(n309), .Y(n543));
sg13g2_nand2_2 U322 (.A(data_o_27_), .B(n304), .Y(n309));
sg13g2_o21ai_1 U323 (.A1(n310), .A2(n304), .B1(n311), .Y(n544));
sg13g2_nand2_2 U324 (.A(data_o_28_), .B(n304), .Y(n311));
sg13g2_o21ai_1 U325 (.A1(n312), .A2(n304), .B1(n313), .Y(n545));
sg13g2_nand2_2 U326 (.A(data_o_29_), .B(n304), .Y(n313));
sg13g2_o21ai_1 U327 (.A1(n314), .A2(n304), .B1(n315), .Y(n546));
sg13g2_nand2_2 U328 (.A(data_o_30_), .B(n304), .Y(n315));
sg13g2_o21ai_1 U329 (.A1(n99), .A2(n203), .B1(n210), .Y(n511));
sg13g2_o21ai_1 U330 (.A1(n168), .A2(n45), .B1(n169), .Y(n501));
sg13g2_o21ai_1 U331 (.A1(n318), .A2(n304), .B1(n319), .Y(n548));
sg13g2_nand2_2 U332 (.A(data_o_24_), .B(n304), .Y(n319));
sg13g2_nand2_2 U333 (.A(n320), .B(n224), .Y(n304));
sg13g2_nor2_2 U334 (.A(n791), .B(n590), .Y(n224));
sg13g2_o21ai_1 U335 (.A1(n303), .A2(n323), .B1(n324), .Y(n549));
sg13g2_nand2_2 U336 (.A(data_o_57_), .B(n323), .Y(n324));
sg13g2_o21ai_1 U337 (.A1(n306), .A2(n323), .B1(n325), .Y(n550));
sg13g2_nand2_2 U338 (.A(data_o_58_), .B(n323), .Y(n325));
sg13g2_o21ai_1 U339 (.A1(n308), .A2(n323), .B1(n326), .Y(n551));
sg13g2_nand2_2 U340 (.A(data_o_59_), .B(n323), .Y(n326));
sg13g2_o21ai_1 U341 (.A1(n310), .A2(n323), .B1(n327), .Y(n552));
sg13g2_nand2_2 U342 (.A(data_o_60_), .B(n323), .Y(n327));
sg13g2_o21ai_1 U343 (.A1(n312), .A2(n323), .B1(n328), .Y(n553));
sg13g2_nand2_2 U344 (.A(data_o_61_), .B(n323), .Y(n328));
sg13g2_o21ai_1 U345 (.A1(n314), .A2(n323), .B1(n329), .Y(n554));
sg13g2_nand2_2 U346 (.A(data_o_62_), .B(n323), .Y(n329));
sg13g2_o21ai_1 U347 (.A1(n316), .A2(n323), .B1(n330), .Y(n555));
sg13g2_nand2_2 U348 (.A(data_o_63_), .B(n323), .Y(n330));
sg13g2_o21ai_1 U349 (.A1(n318), .A2(n323), .B1(n331), .Y(n556));
sg13g2_nand2_2 U350 (.A(data_o_56_), .B(n323), .Y(n331));
sg13g2_nand2_2 U351 (.A(n320), .B(n126), .Y(n323));
sg13g2_nor2_2 U352 (.A(n791), .B(N32), .Y(n126));
sg13g2_inv_4 U353 (.A(N131), .Y(n17));
sg13g2_o21ai_1 U354 (.A1(n303), .A2(n332), .B1(n333), .Y(n557));
sg13g2_nand2_2 U355 (.A(data_o_89_), .B(n332), .Y(n333));
sg13g2_o21ai_1 U356 (.A1(n306), .A2(n332), .B1(n334), .Y(n558));
sg13g2_nand2_2 U357 (.A(data_o_90_), .B(n332), .Y(n334));
sg13g2_o21ai_1 U358 (.A1(n308), .A2(n332), .B1(n335), .Y(n559));
sg13g2_nand2_2 U359 (.A(data_o_91_), .B(n332), .Y(n335));
sg13g2_o21ai_1 U360 (.A1(n310), .A2(n332), .B1(n336), .Y(n560));
sg13g2_nand2_2 U361 (.A(data_o_92_), .B(n332), .Y(n336));
sg13g2_o21ai_1 U362 (.A1(n312), .A2(n332), .B1(n337), .Y(n561));
sg13g2_nand2_2 U363 (.A(data_o_93_), .B(n332), .Y(n337));
sg13g2_o21ai_1 U364 (.A1(n314), .A2(n332), .B1(n338), .Y(n562));
sg13g2_nand2_2 U365 (.A(data_o_94_), .B(n332), .Y(n338));
sg13g2_o21ai_1 U366 (.A1(n316), .A2(n332), .B1(n339), .Y(n563));
sg13g2_nand2_2 U367 (.A(data_o_95_), .B(n332), .Y(n339));
sg13g2_o21ai_1 U368 (.A1(n318), .A2(n332), .B1(n340), .Y(n564));
sg13g2_nand2_2 U369 (.A(data_o_88_), .B(n332), .Y(n340));
sg13g2_nand2_2 U370 (.A(n320), .B(n82), .Y(n332));
sg13g2_nor2_2 U371 (.A(n599), .B(n342), .Y(n320));
sg13g2_o21ai_1 U372 (.A1(n303), .A2(n343), .B1(n344), .Y(n565));
sg13g2_nand2_2 U373 (.A(data_o_121_), .B(n343), .Y(n344));
sg13g2_inv_4 U374 (.A(sbox_data_i_1_), .Y(n303));
sg13g2_o21ai_1 U375 (.A1(n306), .A2(n343), .B1(n345), .Y(n566));
sg13g2_nand2_2 U376 (.A(data_o_122_), .B(n343), .Y(n345));
sg13g2_inv_4 U377 (.A(sbox_data_i_2_), .Y(n306));
sg13g2_o21ai_1 U378 (.A1(n308), .A2(n343), .B1(n346), .Y(n567));
sg13g2_nand2_2 U379 (.A(data_o_123_), .B(n343), .Y(n346));
sg13g2_inv_4 U380 (.A(sbox_data_i_3_), .Y(n308));
sg13g2_o21ai_1 U381 (.A1(n310), .A2(n343), .B1(n347), .Y(n568));
sg13g2_nand2_2 U382 (.A(data_o_124_), .B(n343), .Y(n347));
sg13g2_inv_4 U383 (.A(sbox_data_i_4_), .Y(n310));
sg13g2_o21ai_1 U384 (.A1(n312), .A2(n343), .B1(n348), .Y(n569));
sg13g2_nand2_2 U385 (.A(data_o_125_), .B(n343), .Y(n348));
sg13g2_inv_4 U386 (.A(sbox_data_i_5_), .Y(n312));
sg13g2_o21ai_1 U387 (.A1(n314), .A2(n343), .B1(n349), .Y(n570));
sg13g2_nand2_2 U388 (.A(data_o_126_), .B(n343), .Y(n349));
sg13g2_inv_4 U389 (.A(sbox_data_i_6_), .Y(n314));
sg13g2_o21ai_1 U390 (.A1(n316), .A2(n343), .B1(n350), .Y(n571));
sg13g2_nand2_2 U391 (.A(data_o_127_), .B(n343), .Y(n350));
sg13g2_inv_4 U392 (.A(sbox_data_i_7_), .Y(n316));
sg13g2_o21ai_1 U393 (.A1(n318), .A2(n343), .B1(n351), .Y(n572));
sg13g2_nand2_2 U394 (.A(data_o_120_), .B(n343), .Y(n351));
sg13g2_nand3_1 U395 (.A(n352), .B(n353), .C(n354), .Y(n343));
sg13g2_inv_4 U396 (.A(sbox_data_i_0_), .Y(n318));
sg13g2_nor2_2 U397 (.A(n1), .B(n355), .Y(n573));
sg13g2_inv_4 U398 (.A(N293), .Y(n355));
sg13g2_nor2_2 U399 (.A(n1), .B(n356), .Y(n574));
sg13g2_inv_4 U400 (.A(N294), .Y(n356));
sg13g2_nor2_2 U401 (.A(n1), .B(n357), .Y(n575));
sg13g2_inv_4 U402 (.A(N295), .Y(n357));
sg13g2_nor2_2 U403 (.A(n1), .B(n358), .Y(n576));
sg13g2_inv_4 U404 (.A(N296), .Y(n358));
sg13g2_o21ai_1 U405 (.A1(n20), .A2(n19), .B1(n359), .Y(n577));
sg13g2_nand2_2 U406 (.A(n599), .B(n354), .Y(n359));
sg13g2_inv_4 U407 (.A(n1), .Y(n354));
sg13g2_nand4_1 U408 (.A(n615), .B(n614), .C(n613), .D(n612), .Y(n616));
sg13g2_nand4_1 U409 (.A(n764), .B(n763), .C(n762), .D(n761), .Y(n765));
sg13g2_nand3_1 U410 (.A(n353), .B(n599), .C(n352), .Y(n20));
sg13g2_nand2b_1 U411 (.A_N(data_i_107_), .B(n795), .Y(n807));
sg13g2_a21oi_2 U412 (.A1(n362), .A2(sbox_data_i_7_), .B1(n363), .Y(n361));
sg13g2_nor2_2 U413 (.A(n364), .B(n365), .Y(n363));
sg13g2_nand2_2 U414 (.A(data_o_87_), .B(n29), .Y(n360));
sg13g2_or2_1 U415 (.A(n752), .B(data_i_99_), .X(n808));
sg13g2_nand2b_1 U416 (.A_N(data_i_106_), .B(n795), .Y(n321));
sg13g2_a21oi_2 U417 (.A1(n362), .A2(sbox_data_i_6_), .B1(n368), .Y(n367));
sg13g2_nor2_2 U418 (.A(n369), .B(n365), .Y(n368));
sg13g2_nand2_2 U419 (.A(data_o_86_), .B(n29), .Y(n366));
sg13g2_or2_1 U420 (.A(n752), .B(data_i_98_), .X(n819));
sg13g2_nand2b_1 U421 (.A_N(data_i_105_), .B(n795), .Y(n816));
sg13g2_a21oi_2 U422 (.A1(n362), .A2(sbox_data_i_5_), .B1(n372), .Y(n371));
sg13g2_nor2_2 U423 (.A(n373), .B(n365), .Y(n372));
sg13g2_nand2_2 U424 (.A(data_o_85_), .B(n29), .Y(n370));
sg13g2_or2_1 U425 (.A(n752), .B(data_i_97_), .X(n817));
sg13g2_nand2b_1 U426 (.A_N(data_i_104_), .B(n795), .Y(n810));
sg13g2_a21oi_2 U427 (.A1(n362), .A2(sbox_data_i_4_), .B1(n376), .Y(n375));
sg13g2_nor2_2 U428 (.A(n377), .B(n365), .Y(n376));
sg13g2_nand2_2 U429 (.A(data_o_84_), .B(n29), .Y(n374));
sg13g2_or2_1 U430 (.A(n752), .B(data_i_96_), .X(n809));
sg13g2_nand2_1 U431 (.A(data_o_96_), .B(n868), .Y(n832));
sg13g2_a21oi_2 U432 (.A1(n362), .A2(sbox_data_i_3_), .B1(n380), .Y(n379));
sg13g2_nor2_2 U433 (.A(n22), .B(n365), .Y(n380));
sg13g2_nand2_1 U434 (.A(data_o_97_), .B(n868), .Y(n833));
sg13g2_nand2_2 U435 (.A(n29), .B(data_o_83_), .Y(n378));
sg13g2_nand2_1 U436 (.A(data_o_98_), .B(n868), .Y(n834));
sg13g2_nand2_1 U437 (.A(data_o_99_), .B(n868), .Y(n835));
sg13g2_a21oi_2 U438 (.A1(n362), .A2(sbox_data_i_2_), .B1(n383), .Y(n382));
sg13g2_nor2_2 U439 (.A(n30), .B(n365), .Y(n383));
sg13g2_nand2_1 U440 (.A(data_o_100_), .B(n868), .Y(n836));
sg13g2_nand2_2 U441 (.A(data_o_82_), .B(n29), .Y(n381));
sg13g2_nand2_1 U442 (.A(data_o_101_), .B(n868), .Y(n837));
sg13g2_nand2_1 U443 (.A(data_o_102_), .B(n868), .Y(n838));
sg13g2_a21oi_2 U444 (.A1(n362), .A2(sbox_data_i_1_), .B1(n386), .Y(n385));
sg13g2_nor2_2 U445 (.A(n35), .B(n365), .Y(n386));
sg13g2_nand2_1 U446 (.A(data_o_103_), .B(n868), .Y(n839));
sg13g2_nand2_2 U447 (.A(data_o_81_), .B(n29), .Y(n384));
sg13g2_nand2_1 U448 (.A(data_o_48_), .B(n868), .Y(n840));
sg13g2_nand2_1 U449 (.A(data_o_49_), .B(n868), .Y(n841));
sg13g2_a21oi_2 U450 (.A1(n362), .A2(sbox_data_i_0_), .B1(n389), .Y(n388));
sg13g2_nor2_2 U451 (.A(n40), .B(n365), .Y(n389));
sg13g2_nand2_2 U452 (.A(n390), .B(n587), .Y(n365));
sg13g2_nand2_1 U453 (.A(data_o_50_), .B(n868), .Y(n842));
sg13g2_inv_4 U454 (.A(n390), .Y(n362));
sg13g2_nand2_2 U455 (.A(n167), .B(n352), .Y(n390));
sg13g2_nand2_2 U456 (.A(data_o_80_), .B(n29), .Y(n387));
sg13g2_nand2_1 U457 (.A(data_o_51_), .B(n868), .Y(n843));
sg13g2_nand4_1 U458 (.A(n711), .B(n713), .C(n712), .D(n714), .Y(n715));
sg13g2_a21oi_2 U459 (.A1(n392), .A2(sbox_data_i_7_), .B1(n393), .Y(n391));
sg13g2_nor2_2 U460 (.A(n168), .B(n394), .Y(n393));
sg13g2_nand2_1 U461 (.A(data_o_52_), .B(n868), .Y(n844));
sg13g2_nand2_1 U462 (.A(data_o_53_), .B(n868), .Y(n845));
sg13g2_o21ai_1 U463 (.A1(n587), .A2(n177), .B1(n395), .Y(n454));
sg13g2_a21oi_2 U464 (.A1(n392), .A2(sbox_data_i_6_), .B1(n396), .Y(n395));
sg13g2_nor2_2 U465 (.A(n174), .B(n394), .Y(n396));
sg13g2_nand2_1 U466 (.A(data_o_54_), .B(n868), .Y(n846));
sg13g2_nand2_1 U467 (.A(data_o_55_), .B(n868), .Y(n847));
sg13g2_nand4_1 U468 (.A(state_4_), .B(n352), .C(n599), .D(n444), .Y(n45));
sg13g2_a21oi_2 U469 (.A1(n392), .A2(sbox_data_i_5_), .B1(n398), .Y(n397));
sg13g2_nor2_2 U470 (.A(n178), .B(n394), .Y(n398));
sg13g2_nand2_1 U471 (.A(data_o_80_), .B(n868), .Y(n848));
sg13g2_nand2_1 U472 (.A(data_o_81_), .B(n868), .Y(n849));
sg13g2_o21ai_1 U473 (.A1(n587), .A2(n185), .B1(n399), .Y(n456));
sg13g2_a21oi_2 U474 (.A1(n392), .A2(sbox_data_i_4_), .B1(n400), .Y(n399));
sg13g2_nor2_2 U475 (.A(n182), .B(n394), .Y(n400));
sg13g2_nand2_1 U476 (.A(data_o_82_), .B(n868), .Y(n850));
sg13g2_nand2_1 U477 (.A(data_o_83_), .B(n868), .Y(n851));
sg13g2_nand2_1 U478 (.A(data_o_84_), .B(n868), .Y(n852));
sg13g2_a21oi_2 U479 (.A1(n392), .A2(sbox_data_i_3_), .B1(n402), .Y(n401));
sg13g2_nor2_2 U480 (.A(n186), .B(n394), .Y(n402));
sg13g2_nand2_1 U481 (.A(data_o_85_), .B(n868), .Y(n853));
sg13g2_nand2_1 U482 (.A(data_o_86_), .B(n868), .Y(n854));
sg13g2_o21ai_1 U483 (.A1(n587), .A2(n193), .B1(n403), .Y(n458));
sg13g2_a21oi_2 U484 (.A1(n392), .A2(sbox_data_i_2_), .B1(n404), .Y(n403));
sg13g2_nor2_2 U485 (.A(n190), .B(n394), .Y(n404));
sg13g2_nand2_1 U486 (.A(data_o_87_), .B(n868), .Y(n855));
sg13g2_nand2_1 U487 (.A(data_o_32_), .B(n868), .Y(n856));
sg13g2_inv_4 U488 (.A(n203), .Y(n29));
sg13g2_a21oi_2 U489 (.A1(n392), .A2(sbox_data_i_1_), .B1(n406), .Y(n405));
sg13g2_nor2_2 U490 (.A(n194), .B(n394), .Y(n406));
sg13g2_nand2_1 U491 (.A(data_o_33_), .B(n868), .Y(n857));
sg13g2_nand2_1 U492 (.A(data_o_34_), .B(n868), .Y(n858));
sg13g2_o21ai_1 U493 (.A1(n587), .A2(n201), .B1(n407), .Y(n460));
sg13g2_a21oi_2 U494 (.A1(n392), .A2(sbox_data_i_0_), .B1(n408), .Y(n407));
sg13g2_nor2_2 U495 (.A(n198), .B(n394), .Y(n408));
sg13g2_nand2_2 U496 (.A(n409), .B(n587), .Y(n394));
sg13g2_nand2_1 U497 (.A(data_o_35_), .B(n868), .Y(n859));
sg13g2_inv_4 U498 (.A(n409), .Y(n392));
sg13g2_nand2_2 U499 (.A(n81), .B(n352), .Y(n409));
sg13g2_nor2_2 U500 (.A(n599), .B(n410), .Y(n81));
sg13g2_nand2_1 U501 (.A(data_o_36_), .B(n868), .Y(n860));
sg13g2_o21ai_1 U502 (.A1(n21), .A2(n89), .B1(n411), .Y(n461));
sg13g2_a21oi_2 U503 (.A1(sbox_data_i_7_), .A2(n412), .B1(n413), .Y(n411));
sg13g2_nor2_2 U504 (.A(n279), .B(n414), .Y(n413));
sg13g2_nand2_1 U505 (.A(data_o_37_), .B(n868), .Y(n861));
sg13g2_nand2_1 U506 (.A(data_o_38_), .B(n868), .Y(n862));
sg13g2_o21ai_1 U507 (.A1(n21), .A2(n94), .B1(n415), .Y(n462));
sg13g2_a21oi_2 U508 (.A1(sbox_data_i_6_), .A2(n412), .B1(n416), .Y(n415));
sg13g2_nor2_2 U509 (.A(n282), .B(n414), .Y(n416));
sg13g2_nand2_1 U510 (.A(data_o_39_), .B(n868), .Y(n863));
sg13g2_nand2_1 U511 (.A(data_o_112_), .B(n868), .Y(n864));
sg13g2_o21ai_1 U512 (.A1(n21), .A2(n99), .B1(n417), .Y(n463));
sg13g2_a21oi_2 U513 (.A1(sbox_data_i_5_), .A2(n412), .B1(n418), .Y(n417));
sg13g2_nor2_2 U514 (.A(n285), .B(n414), .Y(n418));
sg13g2_nand2_1 U515 (.A(data_o_113_), .B(n868), .Y(n865));
sg13g2_nand2_1 U516 (.A(data_o_114_), .B(n868), .Y(n866));
sg13g2_o21ai_1 U517 (.A1(n21), .A2(n104), .B1(n419), .Y(n464));
sg13g2_a21oi_2 U518 (.A1(sbox_data_i_4_), .A2(n412), .B1(n420), .Y(n419));
sg13g2_nor2_2 U519 (.A(n288), .B(n414), .Y(n420));
sg13g2_nand2_1 U520 (.A(data_o_115_), .B(n868), .Y(n867));
sg13g2_nand2_1 U521 (.A(data_o_116_), .B(n868), .Y(n820));
sg13g2_o21ai_1 U522 (.A1(n21), .A2(n109), .B1(n421), .Y(n465));
sg13g2_a21oi_2 U523 (.A1(sbox_data_i_3_), .A2(n412), .B1(n422), .Y(n421));
sg13g2_nor2_2 U524 (.A(n291), .B(n414), .Y(n422));
sg13g2_nand2_1 U525 (.A(data_o_117_), .B(n868), .Y(n821));
sg13g2_nand2_1 U526 (.A(data_o_118_), .B(n868), .Y(n822));
sg13g2_o21ai_1 U527 (.A1(n21), .A2(n114), .B1(n423), .Y(n466));
sg13g2_a21oi_2 U528 (.A1(sbox_data_i_2_), .A2(n412), .B1(n424), .Y(n423));
sg13g2_nor2_2 U529 (.A(n294), .B(n414), .Y(n424));
sg13g2_nand2_1 U530 (.A(data_o_119_), .B(n868), .Y(n823));
sg13g2_nand2_1 U531 (.A(data_o_16_), .B(n868), .Y(n824));
sg13g2_o21ai_1 U532 (.A1(n21), .A2(n119), .B1(n425), .Y(n467));
sg13g2_a21oi_2 U533 (.A1(sbox_data_i_1_), .A2(n412), .B1(n426), .Y(n425));
sg13g2_nor2_2 U534 (.A(n297), .B(n414), .Y(n426));
sg13g2_nand2_1 U535 (.A(data_o_17_), .B(n868), .Y(n825));
sg13g2_nand2_1 U536 (.A(data_o_18_), .B(n868), .Y(n826));
sg13g2_o21ai_1 U537 (.A1(n21), .A2(n124), .B1(n427), .Y(n468));
sg13g2_a21oi_2 U538 (.A1(sbox_data_i_0_), .A2(n412), .B1(n428), .Y(n427));
sg13g2_nor2_2 U539 (.A(n300), .B(n414), .Y(n428));
sg13g2_nand2_2 U540 (.A(n429), .B(n587), .Y(n414));
sg13g2_nand2_1 U541 (.A(data_o_19_), .B(n868), .Y(n827));
sg13g2_o21ai_1 U542 (.A1(decrypt_i), .A2(n587), .B1(n429), .Y(n412));
sg13g2_nand2_2 U543 (.A(n127), .B(n82), .Y(n429));
sg13g2_nor2_2 U544 (.A(n342), .B(N30), .Y(n127));
sg13g2_inv_4 U545 (.A(n353), .Y(n342));
sg13g2_nor2_2 U546 (.A(state_4_), .B(N31), .Y(n353));
sg13g2_nand2_1 U547 (.A(data_o_20_), .B(n868), .Y(n828));
sg13g2_nand2_1 U548 (.A(data_o_21_), .B(n868), .Y(n829));
sg13g2_a21oi_2 U549 (.A1(sbox_data_i_7_), .A2(n25), .B1(n432), .Y(n431));
sg13g2_nor2_2 U550 (.A(n27), .B(n128), .Y(n432));
sg13g2_nand2_1 U551 (.A(data_o_22_), .B(n868), .Y(n830));
sg13g2_nand2_2 U552 (.A(data_o_55_), .B(n29), .Y(n430));
sg13g2_nand2_1 U553 (.A(data_o_23_), .B(n868), .Y(n831));
sg13g2_a21oi_2 U555 (.A1(sbox_data_i_6_), .A2(n25), .B1(n435), .Y(n434));
sg13g2_nor2_2 U556 (.A(n27), .B(n135), .Y(n435));
sg13g2_nand2_2 U558 (.A(data_o_54_), .B(n29), .Y(n433));
sg13g2_a21oi_2 U561 (.A1(sbox_data_i_5_), .A2(n25), .B1(n438), .Y(n437));
sg13g2_nor2_2 U562 (.A(n27), .B(n140), .Y(n438));
sg13g2_nand2_2 U564 (.A(data_o_53_), .B(n29), .Y(n436));
sg13g2_a21oi_2 U567 (.A1(sbox_data_i_4_), .A2(n25), .B1(n441), .Y(n440));
sg13g2_nor2_2 U568 (.A(n27), .B(n145), .Y(n441));
sg13g2_nand2_2 U570 (.A(n442), .B(n587), .Y(n27));
sg13g2_inv_4 U571 (.A(n442), .Y(n25));
sg13g2_nand2_2 U572 (.A(n82), .B(n167), .Y(n442));
sg13g2_nor2_2 U573 (.A(n410), .B(N30), .Y(n167));
sg13g2_inv_4 U574 (.A(n443), .Y(n410));
sg13g2_nor2_2 U575 (.A(n444), .B(state_4_), .Y(n443));
sg13g2_nor2_2 U576 (.A(n590), .B(N33), .Y(n82));
sg13g2_nand2_2 U578 (.A(data_o_52_), .B(n29), .Y(n439));
sg13g2_nand2_2 U580 (.A(next_ready_o), .B(n223), .Y(n203));
sg13g2_inv_4 U581 (.A(decrypt_i), .Y(n223));
sg13g2_nand2_2 U583 (.A(decrypt_i), .B(next_ready_o), .Y(n21));
sg13g2_inv_4 U584 (.A(n587), .Y(next_ready_o));
sg13g2_o21ai_1 U585 (.A1(n643), .A2(n642), .B1(n641), .Y(N130));
sg13g2_nor2_2 U588 (.A(N33), .B(N32), .Y(n352));
sg13g2_nor2_2 U589 (.A(data_i_19_), .B(n779), .Y(n679));
sg13g2_o21ai_1 U590 (.A1(n792), .A2(data_i_123_), .B1(n791), .Y(n669));
sg13g2_nand2_2 U591 (.A(data_i_123_), .B(n4), .Y(n12));
sg13g2_nor2_2 U592 (.A(n19), .B(n20), .Y(n4));
sg13g2_inv_4 U593 (.A(start_i), .Y(n19));
sg13g2_a21oi_2 U594 (.A1(n86), .A2(sbox_data_i_2_), .B1(n113), .Y(n112));
sg13g2_nor2_2 U595 (.A(n595), .B(N30), .Y(n795));
sg13g2_nor2_2 U596 (.A(data_i_27_), .B(n787), .Y(n683));
sg13g2_nor2_2 U597 (.A(data_i_93_), .B(n787), .Y(n719));
sg13g2_nor2_2 U598 (.A(data_i_92_), .B(n787), .Y(n695));
sg13g2_nand2_2 U599 (.A(n600), .B(n599), .Y(n787));
sg13g2_nand4_1 U600 (.A(n799), .B(n796), .C(n797), .D(n798), .Y(n800));
sg13g2_nor2_2 U602 (.A(data_i_119_), .B(n783), .Y(n784));
sg13g2_nor2_2 U603 (.A(data_i_54_), .B(n783), .Y(n755));
sg13g2_nand2_2 U604 (.A(n596), .B(N30), .Y(n783));
sg13g2_o21ai_1 U605 (.A1(n11), .A2(n1), .B1(n12), .Y(sbox_data_o_3_));
sg13g2_inv_4 U606 (.A(N128), .Y(n11));
sg13g2_nor2_2 U611 (.A(data_i_63_), .B(n792), .Y(n768));
sg13g2_nor2_2 U613 (.A(data_i_95_), .B(n787), .Y(n788));
sg13g2_inv_4 U614 (.A(n776), .Y(n777));
sg13g2_nor2_2 U615 (.A(data_i_83_), .B(n779), .Y(n675));
sg13g2_a21oi_2 U616 (.A1(n790), .A2(n771), .B1(n770), .Y(n772));
sg13g2_a21oi_2 U617 (.A1(n782), .A2(n651), .B1(n650), .Y(n652));
sg13g2_inv_4 U618 (.A(n786), .Y(n752));
sg13g2_nor2_2 U619 (.A(n595), .B(n599), .Y(n786));
sg13g2_a21oi_2 U620 (.A1(n790), .A2(n646), .B1(n645), .Y(n647));
sg13g2_o21ai_1 U621 (.A1(n802), .A2(n801), .B1(n800), .Y(N124));
sg13g2_nor2_2 U623 (.A(data_i_84_), .B(n779), .Y(n699));
sg13g2_nor2_2 U626 (.A(data_i_28_), .B(n787), .Y(n707));
sg13g2_inv_4 U627 (.A(n694), .Y(n322));
sg13g2_nand2_2 U628 (.A(n341), .B(n578), .Y(n579));
sg13g2_nand2_2 U629 (.A(n579), .B(n791), .Y(n694));
sg13g2_inv_4 U630 (.A(n792), .Y(n341));
sg13g2_inv_4 U631 (.A(data_i_124_), .Y(n578));
sg13g2_nand2_2 U632 (.A(n596), .B(n599), .Y(n792));
sg13g2_nor2_2 U633 (.A(data_i_52_), .B(n783), .Y(n705));
sg13g2_o21ai_1 U634 (.A1(n1), .A2(n2), .B1(n3), .Y(sbox_data_o_7_));
sg13g2_inv_4 U635 (.A(N124), .Y(n2));
sg13g2_o21ai_1 U636 (.A1(n1), .A2(n5), .B1(n6), .Y(sbox_data_o_6_));
sg13g2_a21oi_2 U637 (.A1(n786), .A2(n756), .B1(n755), .Y(n763));
sg13g2_o21ai_1 U638 (.A1(n741), .A2(n742), .B1(n740), .Y(N126));
sg13g2_nand4_1 U639 (.A(n739), .B(n738), .C(n737), .D(n736), .Y(n740));
sg13g2_a21oi_2 U640 (.A1(n795), .A2(n735), .B1(n734), .Y(n736));
sg13g2_o21ai_1 U641 (.A1(data_i_61_), .A2(n792), .B1(N33), .Y(n734));
sg13g2_o21ai_1 U642 (.A1(n618), .A2(n617), .B1(n616), .Y(N131));
sg13g2_nor2_2 U644 (.A(data_i_20_), .B(n779), .Y(n703));
sg13g2_inv_4 U645 (.A(data_i_75_), .Y(n671));
sg13g2_inv_4 U647 (.A(N130), .Y(n15));
sg13g2_nor2_2 U648 (.A(data_i_55_), .B(n783), .Y(n770));
sg13g2_nor2_2 U649 (.A(data_i_51_), .B(n783), .Y(n681));
sg13g2_inv_4 U650 (.A(data_i_67_), .Y(n676));
sg13g2_nand2_2 U651 (.A(n580), .B(n581), .Y(n582));
sg13g2_nand2_2 U652 (.A(n582), .B(n775), .Y(n776));
sg13g2_inv_4 U653 (.A(n779), .Y(n580));
sg13g2_inv_4 U654 (.A(data_i_23_), .Y(n581));
sg13g2_nand2_2 U655 (.A(n600), .B(N30), .Y(n779));
sg13g2_nand2_2 U656 (.A(n774), .B(n786), .Y(n775));
sg13g2_inv_4 U658 (.A(data_i_39_), .Y(n774));
sg13g2_o21ai_1 U660 (.A1(data_i_60_), .A2(n792), .B1(N33), .Y(n709));
sg13g2_a21oi_2 U661 (.A1(n790), .A2(n671), .B1(n670), .Y(n672));
sg13g2_nor2_2 U662 (.A(data_i_91_), .B(n787), .Y(n670));
sg13g2_nand4_1 U663 (.A(n690), .B(n689), .C(n688), .D(n687), .Y(n691));
sg13g2_a21oi_2 U664 (.A1(n676), .A2(n782), .B1(n675), .Y(n677));
sg13g2_o21ai_1 U665 (.A1(data_i_59_), .A2(n792), .B1(N33), .Y(n685));
sg13g2_o21ai_1 U666 (.A1(data_i_127_), .A2(n792), .B1(n791), .Y(n793));
sg13g2_inv_4 U667 (.A(N125), .Y(n5));
sg13g2_a21oi_2 U669 (.A1(n782), .A2(n700), .B1(n699), .Y(n701));
sg13g2_o21ai_1 U670 (.A1(data_i_62_), .A2(n792), .B1(N33), .Y(n759));
sg13g2_a21oi_2 U671 (.A1(n795), .A2(n760), .B1(n759), .Y(n761));
sg13g2_a21oi_2 U672 (.A1(n696), .A2(n790), .B1(n695), .Y(n697));
sg13g2_o21ai_1 U673 (.A1(n716), .A2(n717), .B1(n715), .Y(N127));
sg13g2_nor2_2 U674 (.A(n778), .B(data_i_70_), .Y(n583));
sg13g2_nor2_2 U675 (.A(n583), .B(n749), .Y(n750));
sg13g2_nor2_2 U676 (.A(data_i_86_), .B(n779), .Y(n749));
sg13g2_nor2_2 U678 (.A(n584), .B(data_i_78_), .Y(n585));
sg13g2_nor2_2 U679 (.A(n585), .B(n744), .Y(n745));
sg13g2_nor2_2 U680 (.A(data_i_94_), .B(n787), .Y(n744));
sg13g2_nor2_2 U681 (.A(n598), .B(N30), .Y(n790));
sg13g2_nor2_2 U682 (.A(n586), .B(n601), .Y(n602));
sg13g2_nor2_2 U683 (.A(n778), .B(data_i_64_), .Y(n586));
sg13g2_nor2_2 U684 (.A(n599), .B(n598), .Y(n782));
sg13g2_nor2_2 U685 (.A(data_i_80_), .B(n779), .Y(n601));
sg13g2_o21ai_1 U686 (.A1(data_i_56_), .A2(n792), .B1(N33), .Y(n610));
sg13g2_buf_8 U687 (.A(n45), .X(n587));
sg13g2_nand2_2 U688 (.A(n587), .B(n20), .Y(n1));
sg13g2_buf_8 U689 (.A(decrypt_i), .X(sbox_decrypt_o));
sg13g2_o21ai_1 U691 (.A1(n792), .A2(data_i_120_), .B1(n791), .Y(n589));
sg13g2_inv_4 U692 (.A(n589), .Y(n594));
sg13g2_inv_4 U693 (.A(data_i_72_), .Y(n592));
sg13g2_nor2_2 U694 (.A(data_i_88_), .B(n787), .Y(n591));
sg13g2_a21oi_2 U695 (.A1(n790), .A2(n592), .B1(n591), .Y(n593));
sg13g2_nor2_2 U696 (.A(data_i_112_), .B(n783), .Y(n597));
sg13g2_inv_4 U697 (.A(n597), .Y(n603));
sg13g2_inv_4 U698 (.A(data_i_0_), .Y(n605));
sg13g2_nor2_2 U699 (.A(data_i_16_), .B(n779), .Y(n604));
sg13g2_a21oi_2 U700 (.A1(n782), .A2(n605), .B1(n604), .Y(n615));
sg13g2_inv_4 U701 (.A(data_i_32_), .Y(n607));
sg13g2_nor2_2 U702 (.A(data_i_48_), .B(n783), .Y(n606));
sg13g2_a21oi_2 U703 (.A1(n786), .A2(n607), .B1(n606), .Y(n614));
sg13g2_inv_4 U704 (.A(data_i_8_), .Y(n609));
sg13g2_nor2_2 U705 (.A(data_i_24_), .B(n787), .Y(n608));
sg13g2_a21oi_2 U706 (.A1(n790), .A2(n609), .B1(n608), .Y(n613));
sg13g2_inv_4 U707 (.A(data_i_40_), .Y(n611));
sg13g2_a21oi_2 U708 (.A1(n795), .A2(n611), .B1(n610), .Y(n612));
sg13g2_o21ai_1 U709 (.A1(n792), .A2(data_i_121_), .B1(n791), .Y(n619));
sg13g2_inv_4 U710 (.A(n619), .Y(n623));
sg13g2_inv_4 U711 (.A(data_i_73_), .Y(n621));
sg13g2_nor2_2 U712 (.A(data_i_89_), .B(n787), .Y(n620));
sg13g2_a21oi_2 U713 (.A1(n790), .A2(n621), .B1(n620), .Y(n622));
sg13g2_nor2_2 U714 (.A(data_i_113_), .B(n783), .Y(n624));
sg13g2_inv_4 U715 (.A(n624), .Y(n628));
sg13g2_inv_4 U716 (.A(data_i_65_), .Y(n626));
sg13g2_nor2_2 U717 (.A(data_i_81_), .B(n779), .Y(n625));
sg13g2_a21oi_2 U718 (.A1(n782), .A2(n626), .B1(n625), .Y(n627));
sg13g2_inv_4 U719 (.A(data_i_1_), .Y(n630));
sg13g2_nor2_2 U720 (.A(data_i_17_), .B(n779), .Y(n629));
sg13g2_a21oi_2 U721 (.A1(n782), .A2(n630), .B1(n629), .Y(n640));
sg13g2_inv_4 U722 (.A(data_i_33_), .Y(n632));
sg13g2_nor2_2 U723 (.A(data_i_49_), .B(n783), .Y(n631));
sg13g2_a21oi_2 U724 (.A1(n786), .A2(n632), .B1(n631), .Y(n639));
sg13g2_inv_4 U725 (.A(data_i_9_), .Y(n634));
sg13g2_nor2_2 U726 (.A(data_i_25_), .B(n787), .Y(n633));
sg13g2_a21oi_2 U727 (.A1(n790), .A2(n634), .B1(n633), .Y(n638));
sg13g2_inv_4 U728 (.A(data_i_41_), .Y(n636));
sg13g2_o21ai_1 U729 (.A1(data_i_57_), .A2(n792), .B1(N33), .Y(n635));
sg13g2_a21oi_2 U730 (.A1(n795), .A2(n636), .B1(n635), .Y(n637));
sg13g2_nand4_1 U731 (.A(n640), .B(n639), .C(n638), .D(n637), .Y(n641));
sg13g2_o21ai_1 U732 (.A1(n792), .A2(data_i_122_), .B1(n791), .Y(n644));
sg13g2_inv_4 U733 (.A(n644), .Y(n648));
sg13g2_inv_4 U734 (.A(data_i_74_), .Y(n646));
sg13g2_nor2_2 U735 (.A(data_i_90_), .B(n787), .Y(n645));
sg13g2_nor2_2 U737 (.A(data_i_114_), .B(n783), .Y(n649));
sg13g2_inv_4 U738 (.A(n649), .Y(n653));
sg13g2_inv_4 U739 (.A(data_i_66_), .Y(n651));
sg13g2_nor2_2 U740 (.A(data_i_82_), .B(n779), .Y(n650));
sg13g2_inv_4 U741 (.A(data_i_2_), .Y(n655));
sg13g2_nor2_2 U742 (.A(data_i_18_), .B(n779), .Y(n654));
sg13g2_a21oi_2 U743 (.A1(n782), .A2(n655), .B1(n654), .Y(n665));
sg13g2_inv_4 U744 (.A(data_i_34_), .Y(n657));
sg13g2_nor2_2 U745 (.A(data_i_50_), .B(n783), .Y(n656));
sg13g2_a21oi_2 U746 (.A1(n786), .A2(n657), .B1(n656), .Y(n664));
sg13g2_inv_4 U747 (.A(data_i_10_), .Y(n659));
sg13g2_nor2_2 U748 (.A(data_i_26_), .B(n787), .Y(n658));
sg13g2_a21oi_2 U749 (.A1(n790), .A2(n659), .B1(n658), .Y(n663));
sg13g2_inv_4 U750 (.A(data_i_42_), .Y(n661));
sg13g2_o21ai_1 U751 (.A1(data_i_58_), .A2(n792), .B1(N33), .Y(n660));
sg13g2_a21oi_2 U752 (.A1(n795), .A2(n661), .B1(n660), .Y(n662));
sg13g2_nand4_1 U753 (.A(n665), .B(n664), .C(n663), .D(n662), .Y(n666));
sg13g2_o21ai_1 U754 (.A1(n668), .A2(n667), .B1(n666), .Y(N129));
sg13g2_inv_4 U755 (.A(n669), .Y(n673));
sg13g2_nor2_2 U756 (.A(data_i_115_), .B(n783), .Y(n674));
sg13g2_inv_4 U757 (.A(n674), .Y(n678));
sg13g2_inv_4 U758 (.A(data_i_3_), .Y(n680));
sg13g2_a21oi_2 U759 (.A1(n782), .A2(n680), .B1(n679), .Y(n690));
sg13g2_inv_4 U760 (.A(data_i_35_), .Y(n682));
sg13g2_a21oi_2 U761 (.A1(n786), .A2(n682), .B1(n681), .Y(n689));
sg13g2_inv_4 U762 (.A(data_i_11_), .Y(n684));
sg13g2_a21oi_2 U763 (.A1(n790), .A2(n684), .B1(n683), .Y(n688));
sg13g2_inv_4 U764 (.A(data_i_43_), .Y(n686));
sg13g2_a21oi_2 U765 (.A1(n795), .A2(n686), .B1(n685), .Y(n687));
sg13g2_inv_4 U766 (.A(data_i_76_), .Y(n696));
sg13g2_nor2_2 U767 (.A(data_i_116_), .B(n783), .Y(n698));
sg13g2_inv_4 U768 (.A(n698), .Y(n702));
sg13g2_inv_4 U769 (.A(data_i_68_), .Y(n700));
sg13g2_inv_4 U770 (.A(data_i_4_), .Y(n704));
sg13g2_a21oi_2 U771 (.A1(n782), .A2(n704), .B1(n703), .Y(n714));
sg13g2_inv_4 U772 (.A(data_i_36_), .Y(n706));
sg13g2_a21oi_2 U773 (.A1(n786), .A2(n706), .B1(n705), .Y(n713));
sg13g2_inv_4 U774 (.A(data_i_12_), .Y(n708));
sg13g2_a21oi_2 U775 (.A1(n790), .A2(n708), .B1(n707), .Y(n712));
sg13g2_inv_4 U776 (.A(data_i_44_), .Y(n710));
sg13g2_a21oi_2 U777 (.A1(n795), .A2(n710), .B1(n709), .Y(n711));
sg13g2_o21ai_1 U778 (.A1(n792), .A2(data_i_125_), .B1(n791), .Y(n718));
sg13g2_inv_4 U779 (.A(n718), .Y(n722));
sg13g2_inv_4 U780 (.A(data_i_77_), .Y(n720));
sg13g2_a21oi_2 U781 (.A1(n790), .A2(n720), .B1(n719), .Y(n721));
sg13g2_nor2_2 U782 (.A(data_i_117_), .B(n783), .Y(n723));
sg13g2_inv_4 U783 (.A(n723), .Y(n727));
sg13g2_inv_4 U784 (.A(data_i_69_), .Y(n725));
sg13g2_nor2_2 U785 (.A(data_i_85_), .B(n779), .Y(n724));
sg13g2_a21oi_2 U786 (.A1(n782), .A2(n725), .B1(n724), .Y(n726));
sg13g2_inv_4 U788 (.A(data_i_5_), .Y(n729));
sg13g2_nor2_2 U789 (.A(data_i_21_), .B(n779), .Y(n728));
sg13g2_a21oi_2 U790 (.A1(n782), .A2(n729), .B1(n728), .Y(n739));
sg13g2_inv_4 U791 (.A(data_i_37_), .Y(n731));
sg13g2_nor2_2 U792 (.A(data_i_53_), .B(n783), .Y(n730));
sg13g2_a21oi_2 U793 (.A1(n786), .A2(n731), .B1(n730), .Y(n738));
sg13g2_inv_4 U794 (.A(data_i_13_), .Y(n733));
sg13g2_nor2_2 U795 (.A(data_i_29_), .B(n787), .Y(n732));
sg13g2_a21oi_2 U796 (.A1(n790), .A2(n733), .B1(n732), .Y(n737));
sg13g2_inv_4 U797 (.A(data_i_45_), .Y(n735));
sg13g2_o21ai_1 U798 (.A1(n792), .A2(data_i_126_), .B1(n791), .Y(n743));
sg13g2_inv_4 U799 (.A(n743), .Y(n746));
sg13g2_nor2_2 U800 (.A(data_i_118_), .B(n783), .Y(n748));
sg13g2_inv_4 U801 (.A(n748), .Y(n751));
sg13g2_inv_4 U802 (.A(data_i_6_), .Y(n754));
sg13g2_nor2_2 U803 (.A(data_i_22_), .B(n779), .Y(n753));
sg13g2_a21oi_2 U804 (.A1(n782), .A2(n754), .B1(n753), .Y(n764));
sg13g2_inv_4 U805 (.A(data_i_38_), .Y(n756));
sg13g2_inv_4 U806 (.A(data_i_14_), .Y(n758));
sg13g2_nor2_2 U807 (.A(data_i_30_), .B(n787), .Y(n757));
sg13g2_a21oi_2 U808 (.A1(n790), .A2(n758), .B1(n757), .Y(n762));
sg13g2_inv_4 U809 (.A(data_i_46_), .Y(n760));
sg13g2_inv_4 U810 (.A(data_i_47_), .Y(n769));
sg13g2_a21oi_2 U811 (.A1(n795), .A2(n769), .B1(n768), .Y(n773));
sg13g2_inv_4 U812 (.A(data_i_15_), .Y(n771));
sg13g2_inv_4 U813 (.A(n782), .Y(n778));
sg13g2_inv_4 U814 (.A(data_i_71_), .Y(n781));
sg13g2_nor2_2 U815 (.A(data_i_87_), .B(n779), .Y(n780));
sg13g2_a21oi_2 U816 (.A1(n782), .A2(n781), .B1(n780), .Y(n799));
sg13g2_inv_4 U817 (.A(data_i_103_), .Y(n785));
sg13g2_a21oi_2 U818 (.A1(n786), .A2(n785), .B1(n784), .Y(n798));
sg13g2_inv_4 U819 (.A(data_i_79_), .Y(n789));
sg13g2_a21oi_2 U820 (.A1(n790), .A2(n789), .B1(n788), .Y(n797));
sg13g2_inv_4 U821 (.A(data_i_111_), .Y(n794));
sg13g2_xnor2_1 U822 (.A(N31), .B(n599), .Y(N293));
sg13g2_nand2_2 U823 (.A(N31), .B(N30), .Y(n803));
sg13g2_xnor2_1 U824 (.A(n803), .B(N32), .Y(N294));
sg13g2_nand3_1 U825 (.A(N31), .B(N30), .C(N32), .Y(n804));
sg13g2_xnor2_1 U826 (.A(n804), .B(N33), .Y(N295));
sg13g2_inv_4 U827 (.A(n804), .Y(n805));
sg13g2_nand2_2 U828 (.A(N33), .B(n805), .Y(n806));
sg13g2_xnor2_1 U829 (.A(n806), .B(state_4_), .Y(N296));
sg13g2_dfrbp_1 data_reg_reg_0_ (.CLK(clk), .D(n540), .Q(data_o_0_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_1_ (.CLK(clk), .D(n539), .Q(data_o_1_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_2_ (.CLK(clk), .D(n538), .Q(data_o_2_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_3_ (.CLK(clk), .D(n537), .Q(data_o_3_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_4_ (.CLK(clk), .D(n536), .Q(data_o_4_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_5_ (.CLK(clk), .D(n535), .Q(data_o_5_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_6_ (.CLK(clk), .D(n534), .Q(data_o_6_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_7_ (.CLK(clk), .D(n533), .Q(data_o_7_), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_8_ (.CLK(clk), .D(n532), .Q(data_o_8_), .Q_N(n76), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_9_ (.CLK(clk), .D(n531), .Q(data_o_9_), .Q_N(n72), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_10_ (.CLK(clk), .D(n530), .Q(data_o_10_), .Q_N(n68), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_11_ (.CLK(clk), .D(n529), .Q(data_o_11_), .Q_N(n64), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_12_ (.CLK(clk), .D(n528), .Q(data_o_12_), .Q_N(n60), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_13_ (.CLK(clk), .D(n527), .Q(data_o_13_), .Q_N(n56), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_14_ (.CLK(clk), .D(n526), .Q(data_o_14_), .Q_N(n52), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_15_ (.CLK(clk), .D(n525), .Q(data_o_15_), .Q_N(n46), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_16_ (.CLK(clk), .D(n524), .Q(data_o_16_), .Q_N(n258), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_17_ (.CLK(clk), .D(n523), .Q(data_o_17_), .Q_N(n254), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_18_ (.CLK(clk), .D(n522), .Q(data_o_18_), .Q_N(n250), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_19_ (.CLK(clk), .D(n521), .Q(data_o_19_), .Q_N(n246), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_20_ (.CLK(clk), .D(n520), .Q(data_o_20_), .Q_N(n242), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_21_ (.CLK(clk), .D(n519), .Q(data_o_21_), .Q_N(n238), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_22_ (.CLK(clk), .D(n518), .Q(data_o_22_), .Q_N(n234), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_23_ (.CLK(clk), .D(n517), .Q(data_o_23_), .Q_N(n229), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_24_ (.CLK(clk), .D(n548), .Q(data_o_24_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_25_ (.CLK(clk), .D(n541), .Q(data_o_25_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_26_ (.CLK(clk), .D(n542), .Q(data_o_26_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_27_ (.CLK(clk), .D(n543), .Q(data_o_27_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_28_ (.CLK(clk), .D(n544), .Q(data_o_28_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_29_ (.CLK(clk), .D(n545), .Q(data_o_29_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_30_ (.CLK(clk), .D(n546), .Q(data_o_30_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_31_ (.CLK(clk), .D(n547), .Q(data_o_31_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_32_ (.CLK(clk), .D(n516), .Q(data_o_32_), .Q_N(n120), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_33_ (.CLK(clk), .D(n515), .Q(data_o_33_), .Q_N(n115), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_34_ (.CLK(clk), .D(n514), .Q(data_o_34_), .Q_N(n110), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_35_ (.CLK(clk), .D(n513), .Q(data_o_35_), .Q_N(n105), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_36_ (.CLK(clk), .D(n512), .Q(data_o_36_), .Q_N(n100), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_37_ (.CLK(clk), .D(n511), .Q(data_o_37_), .Q_N(n95), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_38_ (.CLK(clk), .D(n510), .Q(data_o_38_), .Q_N(n90), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_39_ (.CLK(clk), .D(n509), .Q(data_o_39_), .Q_N(n83), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_40_ (.CLK(clk), .D(n508), .Q(data_o_40_), .Q_N(n201), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_41_ (.CLK(clk), .D(n507), .Q(data_o_41_), .Q_N(n197), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_42_ (.CLK(clk), .D(n506), .Q(data_o_42_), .Q_N(n193), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_43_ (.CLK(clk), .D(n505), .Q(data_o_43_), .Q_N(n189), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_44_ (.CLK(clk), .D(n504), .Q(data_o_44_), .Q_N(n185), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_45_ (.CLK(clk), .D(n503), .Q(data_o_45_), .Q_N(n181), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_46_ (.CLK(clk), .D(n502), .Q(data_o_46_), .Q_N(n177), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_47_ (.CLK(clk), .D(n501), .Q(data_o_47_), .Q_N(n173), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_48_ (.CLK(clk), .D(n500), .Q(data_o_48_), .Q_N(n165), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_49_ (.CLK(clk), .D(n499), .Q(data_o_49_), .Q_N(n161), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_50_ (.CLK(clk), .D(n498), .Q(data_o_50_), .Q_N(n157), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_51_ (.CLK(clk), .D(n497), .Q(data_o_51_), .Q_N(n153), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_52_ (.CLK(clk), .D(n496), .Q(data_o_52_), .Q_N(n149), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_53_ (.CLK(clk), .D(n495), .Q(data_o_53_), .Q_N(n144), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_54_ (.CLK(clk), .D(n494), .Q(data_o_54_), .Q_N(n139), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_55_ (.CLK(clk), .D(n493), .Q(data_o_55_), .Q_N(n134), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_56_ (.CLK(clk), .D(n556), .Q(data_o_56_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_57_ (.CLK(clk), .D(n549), .Q(data_o_57_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_58_ (.CLK(clk), .D(n550), .Q(data_o_58_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_59_ (.CLK(clk), .D(n551), .Q(data_o_59_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_60_ (.CLK(clk), .D(n552), .Q(data_o_60_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_61_ (.CLK(clk), .D(n553), .Q(data_o_61_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_62_ (.CLK(clk), .D(n554), .Q(data_o_62_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_63_ (.CLK(clk), .D(n555), .Q(data_o_63_), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_64_ (.CLK(clk), .D(n492), .Q(data_o_64_), .Q_N(n124), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_65_ (.CLK(clk), .D(n491), .Q(data_o_65_), .Q_N(n119), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_66_ (.CLK(clk), .D(n490), .Q(data_o_66_), .Q_N(n114), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_67_ (.CLK(clk), .D(n489), .Q(data_o_67_), .Q_N(n109), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_68_ (.CLK(clk), .D(n488), .Q(data_o_68_), .Q_N(n104), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_69_ (.CLK(clk), .D(n487), .Q(data_o_69_), .Q_N(n99), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_70_ (.CLK(clk), .D(n486), .Q(data_o_70_), .Q_N(n94), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_71_ (.CLK(clk), .D(n485), .Q(data_o_71_), .Q_N(n89), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_72_ (.CLK(clk), .D(n484), .Q(data_o_72_), .Q_N(n79), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_73_ (.CLK(clk), .D(n483), .Q(data_o_73_), .Q_N(n75), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_74_ (.CLK(clk), .D(n482), .Q(data_o_74_), .Q_N(n71), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_75_ (.CLK(clk), .D(n481), .Q(data_o_75_), .Q_N(n67), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_76_ (.CLK(clk), .D(n480), .Q(data_o_76_), .Q_N(n63), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_77_ (.CLK(clk), .D(n479), .Q(data_o_77_), .Q_N(n59), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_78_ (.CLK(clk), .D(n478), .Q(data_o_78_), .Q_N(n55), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_79_ (.CLK(clk), .D(n477), .Q(data_o_79_), .Q_N(n51), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_80_ (.CLK(clk), .D(n476), .Q(data_o_80_), .Q_N(n44), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_81_ (.CLK(clk), .D(n475), .Q(data_o_81_), .Q_N(n39), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_82_ (.CLK(clk), .D(n474), .Q(data_o_82_), .Q_N(n34), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_83_ (.CLK(clk), .D(n473), .Q(data_o_83_), .Q_N(n28), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_84_ (.CLK(clk), .D(n472), .Q(data_o_84_), .Q_N(n145), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_85_ (.CLK(clk), .D(n471), .Q(data_o_85_), .Q_N(n140), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_86_ (.CLK(clk), .D(n470), .Q(data_o_86_), .Q_N(n135), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_87_ (.CLK(clk), .D(n469), .Q(data_o_87_), .Q_N(n128), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_88_ (.CLK(clk), .D(n564), .Q(data_o_88_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_89_ (.CLK(clk), .D(n557), .Q(data_o_89_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_90_ (.CLK(clk), .D(n558), .Q(data_o_90_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_91_ (.CLK(clk), .D(n559), .Q(data_o_91_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_92_ (.CLK(clk), .D(n560), .Q(data_o_92_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_93_ (.CLK(clk), .D(n561), .Q(data_o_93_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_94_ (.CLK(clk), .D(n562), .Q(data_o_94_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_95_ (.CLK(clk), .D(n563), .Q(data_o_95_), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_96_ (.CLK(clk), .D(n468), .Q(data_o_96_), .Q_N(n300), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_97_ (.CLK(clk), .D(n467), .Q(data_o_97_), .Q_N(n297), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_98_ (.CLK(clk), .D(n466), .Q(data_o_98_), .Q_N(n294), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_99_ (.CLK(clk), .D(n465), .Q(data_o_99_), .Q_N(n291), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_100_ (.CLK(clk), .D(n464), .Q(data_o_100_), .Q_N(n288), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_101_ (.CLK(clk), .D(n463), .Q(data_o_101_), .Q_N(n285), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_102_ (.CLK(clk), .D(n462), .Q(data_o_102_), .Q_N(n282), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_103_ (.CLK(clk), .D(n461), .Q(data_o_103_), .Q_N(n279), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_104_ (.CLK(clk), .D(n460), .Q(data_o_104_), .Q_N(n198), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_105_ (.CLK(clk), .D(n459), .Q(data_o_105_), .Q_N(n194), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_106_ (.CLK(clk), .D(n458), .Q(data_o_106_), .Q_N(n190), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_107_ (.CLK(clk), .D(n457), .Q(data_o_107_), .Q_N(n186), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_108_ (.CLK(clk), .D(n456), .Q(data_o_108_), .Q_N(n182), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_109_ (.CLK(clk), .D(n455), .Q(data_o_109_), .Q_N(n178), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_110_ (.CLK(clk), .D(n454), .Q(data_o_110_), .Q_N(n174), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_111_ (.CLK(clk), .D(n453), .Q(data_o_111_), .Q_N(n168), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_112_ (.CLK(clk), .D(n452), .Q(data_o_112_), .Q_N(n40), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_113_ (.CLK(clk), .D(n451), .Q(data_o_113_), .Q_N(n35), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_114_ (.CLK(clk), .D(n450), .Q(data_o_114_), .Q_N(n30), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_115_ (.CLK(clk), .D(n449), .Q(data_o_115_), .Q_N(n22), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_116_ (.CLK(clk), .D(n448), .Q(data_o_116_), .Q_N(n377), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_117_ (.CLK(clk), .D(n447), .Q(data_o_117_), .Q_N(n373), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_118_ (.CLK(clk), .D(n446), .Q(data_o_118_), .Q_N(n369), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_119_ (.CLK(clk), .D(n445), .Q(data_o_119_), .Q_N(n364), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_120_ (.CLK(clk), .D(n572), .Q(data_o_120_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_121_ (.CLK(clk), .D(n565), .Q(data_o_121_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_122_ (.CLK(clk), .D(n566), .Q(data_o_122_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_123_ (.CLK(clk), .D(n567), .Q(data_o_123_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_124_ (.CLK(clk), .D(n568), .Q(data_o_124_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_125_ (.CLK(clk), .D(n569), .Q(data_o_125_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_126_ (.CLK(clk), .D(n570), .Q(data_o_126_), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_127_ (.CLK(clk), .D(n571), .Q(data_o_127_), .RESET_B(reset));
sg13g2_dfrbp_1 ready_o_reg (.CLK(clk), .D(next_ready_o), .Q(ready_o), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_0_ (.CLK(clk), .D(n577), .Q(N30), .Q_N(n599), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_1_ (.CLK(clk), .D(n573), .Q(N31), .Q_N(n444), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_2_ (.CLK(clk), .D(n574), .Q(N32), .Q_N(n590), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_3_ (.CLK(clk), .D(n575), .Q(N33), .Q_N(n791), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_4_ (.CLK(clk), .D(n576), .Q(state_4_), .RESET_B(reset));
endmodule

module sbox (clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, decrypt_i, reset);
input clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, decrypt_i, reset;
output data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_;

sg13g2_xnor2_1 U3 (.A(n32), .B(net26358), .Y(sum1_alph_t_3_));
sg13g2_xnor2_1 U4 (.A(n3), .B(net27689), .Y(sum1_alph_t_2_));
sg13g2_xnor2_1 U5 (.A(net26507), .B(n335), .Y(sum1_alph_t_1_));
sg13g2_nand2_2 U6 (.A(n318), .B(n317), .Y(next_to_invert_2_));
sg13g2_inv_4 U7 (.A(n14), .Y(ah_3_));
sg13g2_nor2_2 U8 (.A(n9), .B(n14), .Y(net27534));
sg13g2_inv_4 U9 (.A(net27539), .Y(n1));
sg13g2_inv_4 U10 (.A(n1), .Y(n15));
sg13g2_o21ai_1 U11 (.A1(n251), .A2(n285), .B1(n224), .Y(n77));
sg13g2_inv_4 U12 (.A(n303), .Y(n304));
sg13g2_inv_4 U13 (.A(n36), .Y(net27426));
sg13g2_inv_4 U14 (.A(n335), .Y(n310));
sg13g2_inv_4 U15 (.A(n102), .Y(n18));
sg13g2_inv_4 U16 (.A(n18), .Y(n25));
sg13g2_nand2_2 U17 (.A(n296), .B(n297), .Y(n30));
sg13g2_nand2_2 U18 (.A(n344), .B(n343), .Y(next_to_invert_3_));
sg13g2_inv_4 U19 (.A(net26517), .Y(n32));
sg13g2_inv_4 U20 (.A(data_i_1_), .Y(net39477));
sg13g2_nand2_2 U21 (.A(n221), .B(net26034), .Y(n33));
sg13g2_inv_4 U22 (.A(n14), .Y(n252));
sg13g2_xnor2_1 U23 (.A(net26739), .B(n35), .Y(n235));
sg13g2_nand4_1 U24 (.A(net26506), .B(net26505), .C(n334), .D(n333), .Y(n318));
sg13g2_inv_4 U25 (.A(n310), .Y(n40));
sg13g2_nand3_1 U26 (.A(net39445), .B(n254), .C(n255), .Y(n44));
sg13g2_nand2_2 U27 (.A(n320), .B(n319), .Y(n307));
sg13g2_nand2_2 U28 (.A(n289), .B(net26662), .Y(n55));
sg13g2_nand2_2 U29 (.A(n248), .B(n247), .Y(n80));
sg13g2_xnor2_1 U30 (.A(n125), .B(n126), .Y(n118));
sg13g2_nand2_2 U31 (.A(net26034), .B(n85), .Y(n84));
sg13g2_nand2_2 U32 (.A(n67), .B(n68), .Y(n244));
sg13g2_inv_4 U33 (.A(n271), .Y(n113));
sg13g2_xnor2_1 U34 (.A(n172), .B(n173), .Y(n171));
sg13g2_xnor2_1 U35 (.A(n66), .B(n86), .Y(n251));
sg13g2_buf_8 U37 (.A(to_invert_2_), .X(n138));
sg13g2_nand2_2 U38 (.A(to_invert_3_), .B(to_invert_1_), .Y(n207));
sg13g2_nor2_2 U39 (.A(n225), .B(n138), .Y(n136));
sg13g2_inv_4 U40 (.A(data_i_0_), .Y(net26281));
sg13g2_nand2_2 U41 (.A(n139), .B(n182), .Y(n227));
sg13g2_nand2_2 U42 (.A(ah_reg_2_), .B(n128), .Y(n162));
sg13g2_xnor2_1 U43 (.A(n76), .B(n280), .Y(n74));
sg13g2_inv_4 U44 (.A(n3), .Y(n249));
sg13g2_inv_4 U45 (.A(n47), .Y(n263));
sg13g2_xnor2_1 U46 (.A(sum1_alph_t_0_), .B(n269), .Y(n51));
sg13g2_inv_4 U47 (.A(n21), .Y(n31));
sg13g2_nand2_2 U48 (.A(net26034), .B(n213), .Y(n212));
sg13g2_nand2_2 U49 (.A(n124), .B(alph_1_), .Y(n155));
sg13g2_mux2_2 U50 (.A0(net39477), .A1(n209), .S(net44790), .X(n47));
sg13g2_nand2_2 U52 (.A(to_invert_0_), .B(n188), .Y(n199));
sg13g2_nand2_2 U53 (.A(n271), .B(n76), .Y(n273));
sg13g2_nand2_2 U54 (.A(net27670), .B(n240), .Y(n319));
sg13g2_nand2_2 U55 (.A(net44791), .B(n110), .Y(n109));
sg13g2_inv_4 U56 (.A(n139), .Y(n225));
sg13g2_nand2_2 U57 (.A(net26359), .B(net26358), .Y(net26361));
sg13g2_inv_4 U58 (.A(net40475), .Y(net26358));
sg13g2_nand2_2 U59 (.A(n66), .B(net44790), .Y(n65));
sg13g2_nand2_2 U60 (.A(n12), .B(n11), .Y(n341));
sg13g2_nand2_2 U61 (.A(to_invert_1_), .B(to_invert_0_), .Y(n187));
sg13g2_nand2_2 U62 (.A(n272), .B(n273), .Y(n68));
sg13g2_o21ai_1 U63 (.A1(n83), .A2(net26034), .B1(n84), .Y(data_o_4_));
sg13g2_o21ai_1 U64 (.A1(net39319), .A2(n278), .B1(n281), .Y(n28));
sg13g2_nand3_1 U65 (.A(n323), .B(n342), .C(n341), .Y(n325));
sg13g2_xnor2_1 U66 (.A(n171), .B(n170), .Y(n114));
sg13g2_nand3_1 U67 (.A(n272), .B(n243), .C(n273), .Y(n245));
sg13g2_nand2_2 U68 (.A(net26034), .B(n79), .Y(n78));
sg13g2_xnor2_1 U69 (.A(n76), .B(n250), .Y(n79));
sg13g2_nand2_2 U70 (.A(net44791), .B(net26750), .Y(n211));
sg13g2_inv_4 U71 (.A(n211), .Y(n326));
sg13g2_nand2_2 U72 (.A(net39279), .B(net39280), .Y(n283));
sg13g2_xnor2_1 U73 (.A(n86), .B(n279), .Y(n85));
sg13g2_inv_4 U74 (.A(n16), .Y(net39280));
sg13g2_nand2_2 U75 (.A(n22), .B(n23), .Y(n317));
sg13g2_nand2_2 U76 (.A(n124), .B(alph_3_), .Y(n179));
sg13g2_xnor2_1 U77 (.A(n92), .B(n250), .Y(n91));
sg13g2_xnor2_1 U78 (.A(n93), .B(n67), .Y(n92));
sg13g2_nand2_2 U79 (.A(n257), .B(alph_2_), .Y(n258));
sg13g2_nand2_2 U80 (.A(n251), .B(n285), .Y(n224));
sg13g2_nand2_2 U81 (.A(net26034), .B(n203), .Y(n202));
sg13g2_inv_4 U82 (.A(n93), .Y(n81));
sg13g2_nand2_2 U83 (.A(n8), .B(n7), .Y(n343));
sg13g2_xnor2_1 U84 (.A(n97), .B(n98), .Y(n96));
sg13g2_nor2_2 U85 (.A(n99), .B(n100), .Y(n98));
sg13g2_nor2_2 U86 (.A(n102), .B(n101), .Y(n97));
sg13g2_xnor2_1 U87 (.A(n103), .B(n104), .Y(n95));
sg13g2_nand2_2 U88 (.A(ah_reg_2_), .B(n105), .Y(n104));
sg13g2_nor2_2 U89 (.A(n106), .B(n107), .Y(n103));
sg13g2_nand2_2 U90 (.A(n124), .B(ah_reg_3_), .Y(n164));
sg13g2_inv_4 U91 (.A(n67), .Y(n243));
sg13g2_nor2_2 U92 (.A(n219), .B(n242), .Y(net40475));
sg13g2_nor2_2 U93 (.A(n46), .B(n9), .Y(n38));
sg13g2_nand2_2 U94 (.A(net26504), .B(net26503), .Y(net26506));
sg13g2_nand4_1 U95 (.A(n325), .B(n324), .C(n282), .D(n283), .Y(n344));
sg13g2_xnor2_1 U96 (.A(n279), .B(n67), .Y(n108));
sg13g2_inv_4 U97 (.A(n184), .Y(n222));
sg13g2_nand2_2 U98 (.A(net26034), .B(n279), .Y(n117));
sg13g2_inv_4 U99 (.A(n222), .Y(n223));
sg13g2_xnor2_1 U100 (.A(n80), .B(n86), .Y(n83));
sg13g2_o21ai_1 U101 (.A1(n77), .A2(net26034), .B1(n78), .Y(data_o_5_));
sg13g2_o21ai_1 U102 (.A1(n108), .A2(net44791), .B1(n109), .Y(data_o_2_));
sg13g2_nand2_2 U103 (.A(n62), .B(n63), .Y(n308));
sg13g2_xnor2_1 U104 (.A(n120), .B(n121), .Y(n119));
sg13g2_nor2_2 U105 (.A(n122), .B(n123), .Y(n121));
sg13g2_nand2_2 U106 (.A(alph_2_), .B(n124), .Y(n120));
sg13g2_inv_4 U107 (.A(n62), .Y(net26727));
sg13g2_nor2_2 U108 (.A(n25), .B(n127), .Y(n126));
sg13g2_nand2_2 U109 (.A(alph_1_), .B(n128), .Y(n125));
sg13g2_inv_4 U110 (.A(n263), .Y(n264));
sg13g2_xnor2_1 U111 (.A(n131), .B(n132), .Y(n130));
sg13g2_nor2_2 U112 (.A(n133), .B(n123), .Y(n132));
sg13g2_inv_4 U113 (.A(n134), .Y(n123));
sg13g2_nand2_2 U114 (.A(alph_3_), .B(n135), .Y(n131));
sg13g2_xnor2_1 U115 (.A(n136), .B(n137), .Y(n135));
sg13g2_inv_4 U116 (.A(net26242), .Y(n265));
sg13g2_nand2_2 U117 (.A(net27343), .B(net27344), .Y(net26482));
sg13g2_nand2_2 U118 (.A(n225), .B(n226), .Y(n228));
sg13g2_nand2_2 U119 (.A(n227), .B(n228), .Y(n151));
sg13g2_nor2_2 U120 (.A(n127), .B(n106), .Y(n140));
sg13g2_inv_4 U121 (.A(n182), .Y(n226));
sg13g2_nand2_2 U122 (.A(n181), .B(n151), .Y(n231));
sg13g2_xnor2_1 U123 (.A(n288), .B(n94), .Y(n146));
sg13g2_nand2_2 U124 (.A(n229), .B(n230), .Y(n232));
sg13g2_nand2_2 U125 (.A(n231), .B(n232), .Y(n99));
sg13g2_inv_4 U126 (.A(n181), .Y(n229));
sg13g2_inv_4 U127 (.A(n151), .Y(n230));
sg13g2_nand2_2 U128 (.A(n15), .B(n264), .Y(n233));
sg13g2_xnor2_1 U130 (.A(n152), .B(n151), .Y(n142));
sg13g2_nand2_2 U131 (.A(alph_2_), .B(n134), .Y(n149));
sg13g2_xnor2_1 U132 (.A(n154), .B(n153), .Y(n134));
sg13g2_xnor2_1 U133 (.A(n155), .B(n156), .Y(n147));
sg13g2_nor2_2 U134 (.A(n99), .B(n127), .Y(n156));
sg13g2_nand2_2 U136 (.A(net27501), .B(n263), .Y(n234));
sg13g2_nand2_2 U137 (.A(n233), .B(n234), .Y(n3));
sg13g2_inv_4 U138 (.A(net26692), .Y(net26242));
sg13g2_nand2_2 U139 (.A(net25922), .B(n259), .Y(next_to_invert_1_));
sg13g2_xnor2_1 U140 (.A(net26245), .B(n19), .Y(n17));
sg13g2_inv_4 U141 (.A(net27693), .Y(n46));
sg13g2_inv_4 U142 (.A(n256), .Y(n54));
sg13g2_xnor2_1 U144 (.A(n164), .B(n165), .Y(n160));
sg13g2_inv_4 U146 (.A(n53), .Y(n327));
sg13g2_nand2_2 U147 (.A(n41), .B(net39428), .Y(n261));
sg13g2_nand2_2 U148 (.A(n105), .B(ah_reg_3_), .Y(n159));
sg13g2_inv_4 U149 (.A(net39445), .Y(net26487));
sg13g2_nand2_2 U150 (.A(n305), .B(n306), .Y(n203));
sg13g2_nand2_2 U151 (.A(net25863), .B(data_i_2_), .Y(n305));
sg13g2_nand2_2 U152 (.A(ah_reg_1_), .B(n128), .Y(n168));
sg13g2_nand2_2 U153 (.A(net27304), .B(n56), .Y(n295));
sg13g2_nand2_2 U154 (.A(ah_reg_2_), .B(n124), .Y(n166));
sg13g2_nor2_2 U155 (.A(n174), .B(n102), .Y(n173));
sg13g2_nand2_2 U156 (.A(net25862), .B(net27197), .Y(n306));
sg13g2_inv_4 U157 (.A(net25862), .Y(net25863));
sg13g2_xnor2_1 U158 (.A(ah_reg_2_), .B(ah_reg_1_), .Y(n174));
sg13g2_nor2_2 U159 (.A(n106), .B(n100), .Y(n172));
sg13g2_xnor2_1 U160 (.A(ah_reg_3_), .B(ah_reg_0_), .Y(n100));
sg13g2_nand3_1 U161 (.A(ah_0_1), .B(n254), .C(n255), .Y(n256));
sg13g2_nor2_2 U162 (.A(n101), .B(n99), .Y(n176));
sg13g2_xnor2_1 U163 (.A(ah_reg_3_), .B(ah_reg_2_), .Y(n101));
sg13g2_nand2_2 U164 (.A(ah_reg_1_), .B(n105), .Y(n175));
sg13g2_inv_4 U165 (.A(n76), .Y(n69));
sg13g2_xnor2_1 U166 (.A(n179), .B(n180), .Y(n178));
sg13g2_nor2_2 U167 (.A(n99), .B(n143), .Y(n180));
sg13g2_xnor2_1 U169 (.A(n147), .B(n148), .Y(n76));
sg13g2_inv_4 U170 (.A(net26493), .Y(net26401));
sg13g2_xnor2_1 U171 (.A(n74), .B(n73), .Y(n71));
sg13g2_inv_4 U172 (.A(n70), .Y(n271));
sg13g2_inv_4 U173 (.A(n42), .Y(n296));
sg13g2_nor2_2 U174 (.A(n142), .B(n122), .Y(n150));
sg13g2_xnor2_1 U175 (.A(n87), .B(n76), .Y(n66));
sg13g2_nand2_2 U176 (.A(n274), .B(n275), .Y(n277));
sg13g2_inv_4 U177 (.A(n13), .Y(n26));
sg13g2_nand2_2 U178 (.A(ah_0_1), .B(n20), .Y(n19));
sg13g2_nand2_2 U179 (.A(net39319), .B(n278), .Y(n281));
sg13g2_inv_4 U180 (.A(n235), .Y(n34));
sg13g2_nand2_2 U181 (.A(net27343), .B(net27344), .Y(net39452));
sg13g2_nand2_2 U182 (.A(n105), .B(ah_reg_0_), .Y(n165));
sg13g2_xnor2_1 U183 (.A(n194), .B(n195), .Y(n177));
sg13g2_nor2_2 U184 (.A(n25), .B(n133), .Y(n195));
sg13g2_xnor2_1 U186 (.A(n189), .B(n190), .Y(n137));
sg13g2_xnor2_1 U187 (.A(n76), .B(n88), .Y(n89));
sg13g2_nand2_2 U188 (.A(n163), .B(n162), .Y(n238));
sg13g2_nand2_2 U189 (.A(n236), .B(n237), .Y(n239));
sg13g2_nand2_2 U190 (.A(n239), .B(n238), .Y(n161));
sg13g2_nand2_2 U191 (.A(alph_0_), .B(n105), .Y(n194));
sg13g2_inv_4 U192 (.A(n162), .Y(n236));
sg13g2_inv_4 U193 (.A(n163), .Y(n237));
sg13g2_xnor2_1 U194 (.A(n181), .B(n198), .Y(n105));
sg13g2_xnor2_1 U195 (.A(n182), .B(n270), .Y(n186));
sg13g2_xnor2_1 U196 (.A(n186), .B(n137), .Y(n106));
sg13g2_nand2_2 U197 (.A(n283), .B(n282), .Y(n7));
sg13g2_nand2_2 U198 (.A(ah_3_), .B(n340), .Y(n36));
sg13g2_nand2_2 U199 (.A(n290), .B(n291), .Y(n240));
sg13g2_inv_4 U200 (.A(net39452), .Y(net26739));
sg13g2_nor2_2 U201 (.A(n241), .B(n265), .Y(n242));
sg13g2_inv_4 U202 (.A(net44791), .Y(n241));
sg13g2_inv_4 U203 (.A(n220), .Y(n219));
sg13g2_inv_4 U204 (.A(net40475), .Y(net39463));
sg13g2_o21ai_1 U205 (.A1(n64), .A2(net26034), .B1(n65), .Y(data_o_7_));
sg13g2_inv_4 U206 (.A(n60), .Y(n300));
sg13g2_nand2_2 U207 (.A(n244), .B(n245), .Y(n64));
sg13g2_xnor2_1 U208 (.A(n66), .B(n86), .Y(n82));
sg13g2_inv_4 U209 (.A(n6), .Y(n289));
sg13g2_nand2_2 U210 (.A(n70), .B(n94), .Y(n247));
sg13g2_nand2_2 U211 (.A(n246), .B(n271), .Y(n248));
sg13g2_nand2_2 U212 (.A(n248), .B(n247), .Y(n88));
sg13g2_inv_4 U213 (.A(n94), .Y(n246));
sg13g2_nand2_2 U214 (.A(to_invert_0_), .B(to_invert_2_), .Y(n188));
sg13g2_xnor2_1 U215 (.A(n152), .B(n181), .Y(n102));
sg13g2_xnor2_1 U216 (.A(n114), .B(n287), .Y(n250));
sg13g2_inv_4 U217 (.A(n287), .Y(n288));
sg13g2_o21ai_1 U218 (.A1(n71), .A2(net44791), .B1(n72), .Y(data_o_6_));
sg13g2_xnor2_1 U219 (.A(n67), .B(n112), .Y(n73));
sg13g2_nand2_2 U220 (.A(net26756), .B(net26692), .Y(net26759));
sg13g2_nand2_2 U221 (.A(n39), .B(n38), .Y(net26991));
sg13g2_inv_4 U222 (.A(n45), .Y(n337));
sg13g2_nand2_2 U223 (.A(n70), .B(n69), .Y(n272));
sg13g2_a21oi_2 U224 (.A1(net44791), .A2(net26242), .B1(n219), .Y(net27611));
sg13g2_nand2_2 U225 (.A(n37), .B(net27535), .Y(n291));
sg13g2_nand2_2 U226 (.A(net26257), .B(n284), .Y(n334));
sg13g2_nand2_2 U227 (.A(net27345), .B(n21), .Y(n293));
sg13g2_xnor2_1 U228 (.A(n191), .B(n184), .Y(n197));
sg13g2_inv_4 U229 (.A(data_i_2_), .Y(net27197));
sg13g2_xnor2_1 U230 (.A(n96), .B(n95), .Y(n275));
sg13g2_xnor2_1 U231 (.A(n50), .B(n49), .Y(next_to_invert_0_));
sg13g2_nand2_2 U232 (.A(net25924), .B(n34), .Y(net25922));
sg13g2_nand2_2 U233 (.A(n52), .B(n51), .Y(n331));
sg13g2_nand2_2 U234 (.A(net27429), .B(net27428), .Y(n35));
sg13g2_nand3_1 U235 (.A(n30), .B(n298), .C(n252), .Y(n253));
sg13g2_inv_4 U236 (.A(n253), .Y(n12));
sg13g2_nand3_1 U237 (.A(n328), .B(n329), .C(n330), .Y(n332));
sg13g2_inv_4 U238 (.A(n58), .Y(n254));
sg13g2_inv_4 U239 (.A(n326), .Y(n255));
sg13g2_nand3_1 U240 (.A(n235), .B(n260), .C(net26991), .Y(n259));
sg13g2_xnor2_1 U241 (.A(n185), .B(n197), .Y(n154));
sg13g2_inv_4 U242 (.A(n142), .Y(n257));
sg13g2_inv_4 U243 (.A(n258), .Y(n141));
sg13g2_xnor2_1 U244 (.A(n96), .B(n95), .Y(n93));
sg13g2_nand2_2 U245 (.A(n260), .B(net26991), .Y(net25924));
sg13g2_nand2_2 U246 (.A(net26989), .B(net26990), .Y(n260));
sg13g2_inv_4 U247 (.A(n39), .Y(net26990));
sg13g2_inv_4 U248 (.A(n38), .Y(net26989));
sg13g2_nand2_2 U249 (.A(ah_2_), .B(net39452), .Y(n62));
sg13g2_nand2_2 U250 (.A(net27674), .B(net26482), .Y(n16));
sg13g2_nand2_2 U251 (.A(net26575), .B(n261), .Y(n39));
sg13g2_nor2_2 U252 (.A(net26487), .B(n3), .Y(net39428));
sg13g2_nand2_2 U253 (.A(net26487), .B(n36), .Y(net27428));
sg13g2_nand2_2 U254 (.A(net26573), .B(n262), .Y(net26575));
sg13g2_nand2_2 U255 (.A(net39445), .B(n249), .Y(n262));
sg13g2_nand2_2 U256 (.A(net27693), .B(n249), .Y(n11));
sg13g2_nand2_2 U257 (.A(net39445), .B(net27426), .Y(net27429));
sg13g2_inv_4 U258 (.A(n41), .Y(net26573));
sg13g2_inv_4 U259 (.A(n263), .Y(net27670));
sg13g2_nand2_2 U260 (.A(n263), .B(net27341), .Y(net27344));
sg13g2_nand2_2 U261 (.A(net26360), .B(net26361), .Y(net39445));
sg13g2_nand2_2 U262 (.A(n26), .B(ah_1_), .Y(n41));
sg13g2_nand2_2 U263 (.A(ah_2_), .B(n26), .Y(n24));
sg13g2_inv_4 U264 (.A(net27539), .Y(net27501));
sg13g2_nand2_2 U265 (.A(n15), .B(n29), .Y(net27502));
sg13g2_nand2_2 U266 (.A(net27539), .B(net44547), .Y(net44749));
sg13g2_nand2_2 U267 (.A(n47), .B(net25877), .Y(net27343));
sg13g2_nand2_2 U268 (.A(net26360), .B(net26361), .Y(ah_0_1));
sg13g2_nand2_2 U269 (.A(ah_1_), .B(n249), .Y(n27));
sg13g2_nand2_2 U270 (.A(n5), .B(net26245), .Y(net26360));
sg13g2_inv_4 U271 (.A(net39463), .Y(net26245));
sg13g2_nand2_2 U272 (.A(net39463), .B(net26669), .Y(net26671));
sg13g2_inv_4 U273 (.A(n5), .Y(net26359));
sg13g2_inv_4 U274 (.A(net26359), .Y(net39323));
sg13g2_inv_4 U275 (.A(n5), .Y(net27345));
sg13g2_inv_4 U276 (.A(data_i_5_), .Y(net26692));
sg13g2_nand2_2 U277 (.A(net26692), .B(net26693), .Y(net26695));
sg13g2_inv_4 U278 (.A(net44790), .Y(net44791));
sg13g2_inv_4 U279 (.A(n57), .Y(net44790));
sg13g2_inv_4 U280 (.A(decrypt_i), .Y(n57));
sg13g2_xnor2_1 U281 (.A(net27691), .B(net27077), .Y(n5));
sg13g2_inv_4 U282 (.A(n48), .Y(net27077));
sg13g2_inv_4 U283 (.A(net27077), .Y(net27078));
sg13g2_nor2_2 U284 (.A(n215), .B(net27623), .Y(net27691));
sg13g2_o21ai_1 U285 (.A1(net26034), .A2(n265), .B1(n33), .Y(net44547));
sg13g2_nand2_2 U286 (.A(data_i_7_), .B(data_i_5_), .Y(net26758));
sg13g2_nand2_2 U287 (.A(data_i_0_), .B(data_i_5_), .Y(net26694));
sg13g2_inv_4 U288 (.A(n48), .Y(n29));
sg13g2_nor2_2 U289 (.A(n218), .B(net44791), .Y(n217));
sg13g2_a21oi_2 U290 (.A1(net44791), .A2(net26287), .B1(n217), .Y(n48));
sg13g2_xnor2_1 U291 (.A(n210), .B(data_i_1_), .Y(n218));
sg13g2_xnor2_1 U292 (.A(data_i_6_), .B(n201), .Y(n210));
sg13g2_xnor2_1 U293 (.A(n210), .B(net26750), .Y(n209));
sg13g2_inv_4 U294 (.A(data_i_3_), .Y(n201));
sg13g2_inv_4 U295 (.A(n201), .Y(net26638));
sg13g2_xnor2_1 U296 (.A(n214), .B(data_i_1_), .Y(n213));
sg13g2_xnor2_1 U297 (.A(data_i_1_), .B(net40403), .Y(n206));
sg13g2_inv_4 U298 (.A(data_i_6_), .Y(net26495));
sg13g2_xnor2_1 U299 (.A(data_i_4_), .B(data_i_6_), .Y(n214));
sg13g2_inv_4 U300 (.A(net26286), .Y(net26287));
sg13g2_inv_4 U301 (.A(data_i_4_), .Y(net26286));
sg13g2_nor2_2 U302 (.A(n216), .B(net44791), .Y(n215));
sg13g2_nor2_2 U303 (.A(net27623), .B(n215), .Y(net27692));
sg13g2_nand2_2 U304 (.A(n267), .B(n266), .Y(n216));
sg13g2_nand2_2 U305 (.A(n204), .B(net26493), .Y(n266));
sg13g2_inv_4 U306 (.A(net26638), .Y(net26493));
sg13g2_nand2_2 U307 (.A(net26401), .B(net26402), .Y(n267));
sg13g2_inv_4 U308 (.A(n204), .Y(net26402));
sg13g2_nor2_2 U309 (.A(net27621), .B(net26495), .Y(net27623));
sg13g2_xnor2_1 U310 (.A(data_i_7_), .B(data_i_4_), .Y(net40403));
sg13g2_nand2_2 U311 (.A(net26034), .B(n91), .Y(n90));
sg13g2_nand2_2 U312 (.A(to_invert_1_), .B(to_invert_2_), .Y(n192));
sg13g2_xnor2_1 U313 (.A(n207), .B(n192), .Y(n190));
sg13g2_inv_4 U314 (.A(net25877), .Y(net27341));
sg13g2_nor2_2 U315 (.A(n102), .B(n107), .Y(n163));
sg13g2_nand2_2 U316 (.A(net27078), .B(net27501), .Y(n292));
sg13g2_nand2_2 U317 (.A(net27501), .B(net44748), .Y(n268));
sg13g2_nand2_2 U318 (.A(n268), .B(net44749), .Y(n42));
sg13g2_inv_4 U319 (.A(net44547), .Y(net44748));
sg13g2_inv_4 U320 (.A(data_i_0_), .Y(net26693));
sg13g2_o21ai_1 U321 (.A1(net26034), .A2(net40367), .B1(n212), .Y(n200));
sg13g2_nand2_2 U322 (.A(n202), .B(n315), .Y(n269));
sg13g2_inv_4 U323 (.A(n193), .Y(n270));
sg13g2_inv_4 U324 (.A(n6), .Y(n340));
sg13g2_xnor2_1 U325 (.A(n66), .B(n94), .Y(n144));
sg13g2_nand2_2 U326 (.A(ah_0_1), .B(net26482), .Y(n278));
sg13g2_xnor2_1 U327 (.A(n75), .B(n114), .Y(n87));
sg13g2_xnor2_1 U328 (.A(n94), .B(n82), .Y(n116));
sg13g2_inv_4 U329 (.A(net44791), .Y(net26034));
sg13g2_inv_4 U330 (.A(net26281), .Y(net26750));
sg13g2_xnor2_1 U331 (.A(n196), .B(n154), .Y(n152));
sg13g2_inv_4 U332 (.A(net44791), .Y(net27621));
sg13g2_nand2_2 U333 (.A(n75), .B(n81), .Y(n276));
sg13g2_nand2_2 U334 (.A(n276), .B(n277), .Y(n70));
sg13g2_inv_4 U335 (.A(n75), .Y(n274));
sg13g2_nand2_2 U336 (.A(net39323), .B(n31), .Y(net27347));
sg13g2_xnor2_1 U337 (.A(data_i_2_), .B(net40403), .Y(n221));
sg13g2_inv_4 U338 (.A(data_i_7_), .Y(net26756));
sg13g2_buf_8 U339 (.A(net26756), .X(net40367));
sg13g2_nand2_2 U340 (.A(n113), .B(net44791), .Y(n72));
sg13g2_o21ai_1 U341 (.A1(to_invert_3_), .A2(n138), .B1(n223), .Y(n181));
sg13g2_inv_4 U342 (.A(n269), .Y(net26669));
sg13g2_xnor2_1 U343 (.A(n175), .B(n176), .Y(n170));
sg13g2_nand2_2 U344 (.A(n6), .B(net27500), .Y(n290));
sg13g2_inv_4 U345 (.A(net27692), .Y(net27304));
sg13g2_xnor2_1 U346 (.A(n115), .B(n159), .Y(n158));
sg13g2_nand2_2 U347 (.A(to_invert_3_), .B(to_invert_2_), .Y(n184));
sg13g2_inv_4 U348 (.A(n73), .Y(n86));
sg13g2_xnor2_1 U349 (.A(n112), .B(n250), .Y(n111));
sg13g2_xnor2_1 U350 (.A(n118), .B(n119), .Y(n112));
sg13g2_inv_4 U351 (.A(n17), .Y(net39279));
sg13g2_nand2_2 U352 (.A(n17), .B(n16), .Y(n282));
sg13g2_inv_4 U353 (.A(n11), .Y(net25870));
sg13g2_nand2_2 U354 (.A(n304), .B(n309), .Y(n312));
sg13g2_xnor2_1 U355 (.A(n94), .B(n111), .Y(n110));
sg13g2_buf_8 U356 (.A(n87), .X(n279));
sg13g2_inv_4 U357 (.A(n75), .Y(n280));
sg13g2_inv_4 U358 (.A(net25860), .Y(net39319));
sg13g2_inv_4 U359 (.A(n28), .Y(net26504));
sg13g2_nand2_2 U360 (.A(ah_3_), .B(n249), .Y(n63));
sg13g2_inv_4 U361 (.A(n43), .Y(n297));
sg13g2_nand2_2 U362 (.A(n28), .B(n27), .Y(net26505));
sg13g2_nand2_2 U363 (.A(net26506), .B(net26505), .Y(n22));
sg13g2_inv_4 U364 (.A(n27), .Y(net26503));
sg13g2_buf_8 U365 (.A(n29), .X(net25860));
sg13g2_inv_4 U366 (.A(n29), .Y(net27500));
sg13g2_nand2_2 U367 (.A(n221), .B(net26034), .Y(n220));
sg13g2_nand2_2 U368 (.A(net27343), .B(net27344), .Y(n21));
sg13g2_nand2_2 U369 (.A(n55), .B(n313), .Y(net27693));
sg13g2_inv_4 U370 (.A(net26662), .Y(net27689));
sg13g2_nand2_2 U371 (.A(n323), .B(ah_3_), .Y(n284));
sg13g2_inv_4 U372 (.A(n307), .Y(n323));
sg13g2_nand2_2 U373 (.A(n293), .B(net27347), .Y(net27674));
sg13g2_inv_4 U374 (.A(n185), .Y(n183));
sg13g2_inv_4 U375 (.A(n275), .Y(n285));
sg13g2_nor2_2 U376 (.A(net44791), .B(n206), .Y(n286));
sg13g2_inv_4 U377 (.A(net27078), .Y(net27535));
sg13g2_nand2_2 U378 (.A(sum1_alph_t_0_), .B(net27692), .Y(n294));
sg13g2_inv_4 U379 (.A(n115), .Y(n287));
sg13g2_xnor2_1 U380 (.A(n160), .B(n161), .Y(n115));
sg13g2_nand2_2 U381 (.A(n290), .B(n291), .Y(n2));
sg13g2_a21oi_2 U382 (.A1(net44791), .A2(net26713), .B1(n286), .Y(net27539));
sg13g2_nand2_2 U383 (.A(net27502), .B(n292), .Y(n20));
sg13g2_xnor2_1 U384 (.A(n129), .B(n130), .Y(n67));
sg13g2_xnor2_1 U385 (.A(n140), .B(n141), .Y(n129));
sg13g2_o21ai_1 U386 (.A1(net26034), .A2(n89), .B1(n90), .Y(data_o_3_));
sg13g2_nand2_2 U387 (.A(n61), .B(n40), .Y(n311));
sg13g2_inv_4 U388 (.A(n106), .Y(n124));
sg13g2_inv_4 U389 (.A(n4), .Y(net26662));
sg13g2_nor2_2 U390 (.A(n100), .B(n102), .Y(n169));
sg13g2_nand2_2 U391 (.A(net27347), .B(n293), .Y(ah_1_));
sg13g2_o21ai_1 U392 (.A1(net26034), .A2(net40367), .B1(n212), .Y(net25877));
sg13g2_nand2_2 U393 (.A(n295), .B(n294), .Y(n43));
sg13g2_nand2_2 U394 (.A(n43), .B(n42), .Y(n298));
sg13g2_nand2_2 U395 (.A(n296), .B(n297), .Y(n299));
sg13g2_nand2_2 U396 (.A(n299), .B(n298), .Y(n13));
sg13g2_nand2_2 U397 (.A(net27611), .B(n269), .Y(n316));
sg13g2_nand2_2 U398 (.A(n60), .B(data_i_2_), .Y(n301));
sg13g2_nand2_2 U399 (.A(n300), .B(net27197), .Y(n302));
sg13g2_nand2_2 U400 (.A(n301), .B(n302), .Y(n59));
sg13g2_nand2_2 U401 (.A(n342), .B(n341), .Y(n10));
sg13g2_nand2_2 U402 (.A(n253), .B(net25870), .Y(n342));
sg13g2_nand2_2 U403 (.A(n320), .B(n319), .Y(n9));
sg13g2_nand2_2 U404 (.A(n6), .B(n4), .Y(n313));
sg13g2_inv_4 U405 (.A(n340), .Y(n335));
sg13g2_nand2_2 U406 (.A(n308), .B(n310), .Y(n303));
sg13g2_nor2_2 U407 (.A(n187), .B(n193), .Y(n189));
sg13g2_xnor2_1 U408 (.A(n196), .B(n153), .Y(n198));
sg13g2_o21ai_1 U409 (.A1(n192), .A2(n207), .B1(to_invert_1_), .Y(n196));
sg13g2_nand2_2 U410 (.A(to_invert_3_), .B(to_invert_1_), .Y(n191));
sg13g2_nand2_2 U411 (.A(net26034), .B(n146), .Y(n145));
sg13g2_inv_4 U412 (.A(n99), .Y(n128));
sg13g2_xnor2_1 U413 (.A(n168), .B(n169), .Y(n167));
sg13g2_xnor2_1 U414 (.A(n177), .B(n178), .Y(n94));
sg13g2_o21ai_1 U415 (.A1(to_invert_0_), .A2(n192), .B1(n199), .Y(n153));
sg13g2_xnor2_1 U416 (.A(n187), .B(n188), .Y(n182));
sg13g2_nand2_2 U417 (.A(to_invert_0_), .B(to_invert_3_), .Y(n185));
sg13g2_xnor2_1 U418 (.A(n158), .B(n157), .Y(n75));
sg13g2_xnor2_1 U419 (.A(n166), .B(n167), .Y(n157));
sg13g2_inv_4 U420 (.A(n56), .Y(sum1_alph_t_0_));
sg13g2_nand2_2 U421 (.A(net44547), .B(net25877), .Y(n321));
sg13g2_nand2_2 U422 (.A(n54), .B(n53), .Y(n328));
sg13g2_nand2_2 U423 (.A(net27674), .B(n20), .Y(n53));
sg13g2_nand2_2 U424 (.A(net26758), .B(net26759), .Y(n60));
sg13g2_nor2_2 U425 (.A(n58), .B(n326), .Y(n56));
sg13g2_nand2_2 U426 (.A(net26727), .B(net26728), .Y(n309));
sg13g2_nand2_2 U427 (.A(n308), .B(n309), .Y(n61));
sg13g2_inv_4 U428 (.A(n63), .Y(net26728));
sg13g2_buf_8 U429 (.A(data_i_2_), .X(net26713));
sg13g2_nand2_2 U430 (.A(n24), .B(net27534), .Y(n333));
sg13g2_nand2_2 U431 (.A(net26695), .B(net26694), .Y(n204));
sg13g2_nand2_2 U432 (.A(n312), .B(n311), .Y(n49));
sg13g2_inv_4 U433 (.A(n204), .Y(net25862));
sg13g2_nand2_2 U434 (.A(net26662), .B(n289), .Y(n314));
sg13g2_nand2_2 U435 (.A(n313), .B(n314), .Y(ah_2_));
sg13g2_nand2_2 U436 (.A(net26665), .B(net26401), .Y(n315));
sg13g2_inv_4 U437 (.A(net26034), .Y(net26665));
sg13g2_nand2_2 U438 (.A(n316), .B(net26671), .Y(n4));
sg13g2_xnor2_1 U439 (.A(n149), .B(n150), .Y(n148));
sg13g2_nand2_2 U440 (.A(net27611), .B(net27341), .Y(n322));
sg13g2_nand2_2 U441 (.A(n327), .B(n44), .Y(n329));
sg13g2_inv_4 U442 (.A(n37), .Y(n6));
sg13g2_nand2_2 U443 (.A(net26517), .B(net26516), .Y(n320));
sg13g2_inv_4 U444 (.A(net27670), .Y(net26516));
sg13g2_inv_4 U445 (.A(n2), .Y(net26517));
sg13g2_nand2_2 U446 (.A(n307), .B(n10), .Y(n324));
sg13g2_inv_4 U447 (.A(net27345), .Y(net26507));
sg13g2_nand2_2 U448 (.A(n321), .B(n322), .Y(n14));
sg13g2_nand2_2 U449 (.A(n324), .B(n325), .Y(n8));
sg13g2_nand2_2 U450 (.A(n329), .B(n328), .Y(n52));
sg13g2_nand2_2 U451 (.A(n332), .B(n331), .Y(n50));
sg13g2_inv_4 U452 (.A(n51), .Y(n330));
sg13g2_nand2_2 U453 (.A(n334), .B(n333), .Y(n23));
sg13g2_inv_4 U454 (.A(n24), .Y(net26257));
sg13g2_nor2_2 U455 (.A(n59), .B(net44791), .Y(n58));
sg13g2_nand2_2 U456 (.A(n45), .B(n200), .Y(n338));
sg13g2_nand2_2 U457 (.A(n337), .B(n336), .Y(n339));
sg13g2_nand2_2 U458 (.A(n339), .B(n338), .Y(n37));
sg13g2_inv_4 U459 (.A(n200), .Y(n336));
sg13g2_nand2_2 U460 (.A(n223), .B(n183), .Y(n139));
sg13g2_o21ai_1 U461 (.A1(net26034), .A2(n144), .B1(n145), .Y(data_o_0_));
sg13g2_a21oi_2 U462 (.A1(net44791), .A2(net26713), .B1(n205), .Y(n45));
sg13g2_nor2_2 U463 (.A(n206), .B(net44791), .Y(n205));
sg13g2_o21ai_1 U464 (.A1(net26034), .A2(n116), .B1(n117), .Y(data_o_1_));
sg13g2_dfrbp_1 ah_reg_reg_0_ (.CLK(clk), .D(net39445), .Q(ah_reg_0_), .RESET_B(reset));
sg13g2_dfrbp_1 ah_reg_reg_1_ (.CLK(clk), .D(ah_1_), .Q(ah_reg_1_), .Q_N(n107), .RESET_B(reset));
sg13g2_dfrbp_1 ah_reg_reg_2_ (.CLK(clk), .D(ah_2_), .Q(ah_reg_2_), .RESET_B(reset));
sg13g2_dfrbp_1 ah_reg_reg_3_ (.CLK(clk), .D(ah_3_), .Q(ah_reg_3_), .RESET_B(reset));
sg13g2_dfrbp_1 alph_reg_0_ (.CLK(clk), .D(sum1_alph_t_0_), .Q(alph_0_), .Q_N(n127), .RESET_B(reset));
sg13g2_dfrbp_1 alph_reg_1_ (.CLK(clk), .D(sum1_alph_t_1_), .Q(alph_1_), .Q_N(n133), .RESET_B(reset));
sg13g2_dfrbp_1 alph_reg_2_ (.CLK(clk), .D(sum1_alph_t_2_), .Q(alph_2_), .Q_N(n143), .RESET_B(reset));
sg13g2_dfrbp_1 alph_reg_3_ (.CLK(clk), .D(sum1_alph_t_3_), .Q(alph_3_), .Q_N(n122), .RESET_B(reset));
sg13g2_dfrbp_1 to_invert_reg_0_ (.CLK(clk), .D(next_to_invert_0_), .Q(to_invert_0_), .RESET_B(reset));
sg13g2_dfrbp_1 to_invert_reg_1_ (.CLK(clk), .D(next_to_invert_1_), .Q(to_invert_1_), .RESET_B(reset));
sg13g2_dfrbp_1 to_invert_reg_2_ (.CLK(clk), .D(next_to_invert_2_), .Q(to_invert_2_), .RESET_B(reset));
sg13g2_dfrbp_1 to_invert_reg_3_ (.CLK(clk), .D(next_to_invert_3_), .Q(to_invert_3_), .Q_N(n193), .RESET_B(reset));
endmodule

module mixcolum (clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_i_8_, data_i_9_, data_i_10_, data_i_11_, data_i_12_, data_i_13_, data_i_14_, data_i_15_, data_i_16_, data_i_17_, data_i_18_, data_i_19_, data_i_20_, data_i_21_, data_i_22_, data_i_23_, data_i_24_, data_i_25_, data_i_26_, data_i_27_, data_i_28_, data_i_29_, data_i_30_, data_i_31_, data_i_32_, data_i_33_, data_i_34_, data_i_35_, data_i_36_, data_i_37_, data_i_38_, data_i_39_, data_i_40_, data_i_41_, data_i_42_, data_i_43_, data_i_44_, data_i_45_, data_i_46_, data_i_47_, data_i_48_, data_i_49_, data_i_50_, data_i_51_, data_i_52_, data_i_53_, data_i_54_, data_i_55_, data_i_56_, data_i_57_, data_i_58_, data_i_59_, data_i_60_, data_i_61_, data_i_62_, data_i_63_, data_i_64_, data_i_65_, data_i_66_, data_i_67_, data_i_68_, data_i_69_, data_i_70_, data_i_71_, data_i_72_, data_i_73_, data_i_74_, data_i_75_, data_i_76_, data_i_77_, data_i_78_, data_i_79_, data_i_80_, data_i_81_, data_i_82_, data_i_83_, data_i_84_, data_i_85_, data_i_86_, data_i_87_, data_i_88_, data_i_89_, data_i_90_, data_i_91_, data_i_92_, data_i_93_, data_i_94_, data_i_95_, data_i_96_, data_i_97_, data_i_98_, data_i_99_, data_i_100_, data_i_101_, data_i_102_, data_i_103_, data_i_104_, data_i_105_, data_i_106_, data_i_107_, data_i_108_, data_i_109_, data_i_110_, data_i_111_, data_i_112_, data_i_113_, data_i_114_, data_i_115_, data_i_116_, data_i_117_, data_i_118_, data_i_119_, data_i_120_, data_i_121_, data_i_122_, data_i_123_, data_i_124_, data_i_125_, data_i_126_, data_i_127_, data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_, data_o_32_, data_o_33_, data_o_34_, data_o_35_, data_o_36_, data_o_37_, data_o_38_, data_o_39_, data_o_40_, data_o_41_, data_o_42_, data_o_43_, data_o_44_, data_o_45_, data_o_46_, data_o_47_, data_o_48_, data_o_49_, data_o_50_, data_o_51_, data_o_52_, data_o_53_, data_o_54_, data_o_55_, data_o_56_, data_o_57_, data_o_58_, data_o_59_, data_o_60_, data_o_61_, data_o_62_, data_o_63_, data_o_64_, data_o_65_, data_o_66_, data_o_67_, data_o_68_, data_o_69_, data_o_70_, data_o_71_, data_o_72_, data_o_73_, data_o_74_, data_o_75_, data_o_76_, data_o_77_, data_o_78_, data_o_79_, data_o_80_, data_o_81_, data_o_82_, data_o_83_, data_o_84_, data_o_85_, data_o_86_, data_o_87_, data_o_88_, data_o_89_, data_o_90_, data_o_91_, data_o_92_, data_o_93_, data_o_94_, data_o_95_, data_o_96_, data_o_97_, data_o_98_, data_o_99_, data_o_100_, data_o_101_, data_o_102_, data_o_103_, data_o_104_, data_o_105_, data_o_106_, data_o_107_, data_o_108_, data_o_109_, data_o_110_, data_o_111_, data_o_112_, data_o_113_, data_o_114_, data_o_115_, data_o_116_, data_o_117_, data_o_118_, data_o_119_, data_o_120_, data_o_121_, data_o_122_, data_o_123_, data_o_124_, data_o_125_, data_o_126_, data_o_127_, decrypt_i, ready_o, reset, start_i);
input clk, data_i_0_, data_i_1_, data_i_2_, data_i_3_, data_i_4_, data_i_5_, data_i_6_, data_i_7_, data_i_8_, data_i_9_, data_i_10_, data_i_11_, data_i_12_, data_i_13_, data_i_14_, data_i_15_, data_i_16_, data_i_17_, data_i_18_, data_i_19_, data_i_20_, data_i_21_, data_i_22_, data_i_23_, data_i_24_, data_i_25_, data_i_26_, data_i_27_, data_i_28_, data_i_29_, data_i_30_, data_i_31_, data_i_32_, data_i_33_, data_i_34_, data_i_35_, data_i_36_, data_i_37_, data_i_38_, data_i_39_, data_i_40_, data_i_41_, data_i_42_, data_i_43_, data_i_44_, data_i_45_, data_i_46_, data_i_47_, data_i_48_, data_i_49_, data_i_50_, data_i_51_, data_i_52_, data_i_53_, data_i_54_, data_i_55_, data_i_56_, data_i_57_, data_i_58_, data_i_59_, data_i_60_, data_i_61_, data_i_62_, data_i_63_, data_i_64_, data_i_65_, data_i_66_, data_i_67_, data_i_68_, data_i_69_, data_i_70_, data_i_71_, data_i_72_, data_i_73_, data_i_74_, data_i_75_, data_i_76_, data_i_77_, data_i_78_, data_i_79_, data_i_80_, data_i_81_, data_i_82_, data_i_83_, data_i_84_, data_i_85_, data_i_86_, data_i_87_, data_i_88_, data_i_89_, data_i_90_, data_i_91_, data_i_92_, data_i_93_, data_i_94_, data_i_95_, data_i_96_, data_i_97_, data_i_98_, data_i_99_, data_i_100_, data_i_101_, data_i_102_, data_i_103_, data_i_104_, data_i_105_, data_i_106_, data_i_107_, data_i_108_, data_i_109_, data_i_110_, data_i_111_, data_i_112_, data_i_113_, data_i_114_, data_i_115_, data_i_116_, data_i_117_, data_i_118_, data_i_119_, data_i_120_, data_i_121_, data_i_122_, data_i_123_, data_i_124_, data_i_125_, data_i_126_, data_i_127_, decrypt_i, reset, start_i;
output data_o_0_, data_o_1_, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_, data_o_32_, data_o_33_, data_o_34_, data_o_35_, data_o_36_, data_o_37_, data_o_38_, data_o_39_, data_o_40_, data_o_41_, data_o_42_, data_o_43_, data_o_44_, data_o_45_, data_o_46_, data_o_47_, data_o_48_, data_o_49_, data_o_50_, data_o_51_, data_o_52_, data_o_53_, data_o_54_, data_o_55_, data_o_56_, data_o_57_, data_o_58_, data_o_59_, data_o_60_, data_o_61_, data_o_62_, data_o_63_, data_o_64_, data_o_65_, data_o_66_, data_o_67_, data_o_68_, data_o_69_, data_o_70_, data_o_71_, data_o_72_, data_o_73_, data_o_74_, data_o_75_, data_o_76_, data_o_77_, data_o_78_, data_o_79_, data_o_80_, data_o_81_, data_o_82_, data_o_83_, data_o_84_, data_o_85_, data_o_86_, data_o_87_, data_o_88_, data_o_89_, data_o_90_, data_o_91_, data_o_92_, data_o_93_, data_o_94_, data_o_95_, data_o_96_, data_o_97_, data_o_98_, data_o_99_, data_o_100_, data_o_101_, data_o_102_, data_o_103_, data_o_104_, data_o_105_, data_o_106_, data_o_107_, data_o_108_, data_o_109_, data_o_110_, data_o_111_, data_o_112_, data_o_113_, data_o_114_, data_o_115_, data_o_116_, data_o_117_, data_o_118_, data_o_119_, data_o_120_, data_o_121_, data_o_122_, data_o_123_, data_o_124_, data_o_125_, data_o_126_, data_o_127_, ready_o;

sg13g2_nand3_1 U1 (.A(n430), .B(n46), .C(n429), .Y(n789));
sg13g2_nand3_1 U2 (.A(n392), .B(n57), .C(n391), .Y(n770));
sg13g2_o21ai_1 U3 (.A1(n1), .A2(n2), .B1(n3), .Y(n663));
sg13g2_a21oi_2 U4 (.A1(outx_31_), .A2(n4), .B1(n5), .Y(n3));
sg13g2_inv_4 U5 (.A(outy_5_), .Y(n28));
sg13g2_o21ai_1 U6 (.A1(n8), .A2(n9), .B1(n10), .Y(n664));
sg13g2_a21oi_2 U7 (.A1(n11), .A2(outy_31_), .B1(n12), .Y(n10));
sg13g2_nor2_2 U8 (.A(n13), .B(n14), .Y(n12));
sg13g2_o21ai_1 U9 (.A1(n15), .A2(n16), .B1(n17), .Y(n665));
sg13g2_inv_4 U10 (.A(n28), .Y(n35));
sg13g2_nor2_2 U11 (.A(n13), .B(n20), .Y(n19));
sg13g2_inv_4 U12 (.A(outx_31_), .Y(n13));
sg13g2_o21ai_1 U13 (.A1(n1), .A2(n153), .B1(n154), .Y(n702));
sg13g2_o21ai_1 U14 (.A1(n1), .A2(n307), .B1(n308), .Y(n744));
sg13g2_o21ai_1 U15 (.A1(n1), .A2(n32), .B1(n33), .Y(n669));
sg13g2_o21ai_1 U16 (.A1(n8), .A2(n25), .B1(n26), .Y(n667));
sg13g2_a21oi_2 U17 (.A1(outy_30_), .A2(n11), .B1(n27), .Y(n26));
sg13g2_nor2_2 U18 (.A(n14), .B(n902), .Y(n27));
sg13g2_o21ai_1 U19 (.A1(n15), .A2(n29), .B1(n30), .Y(n668));
sg13g2_a21oi_2 U20 (.A1(outy_30_), .A2(n18), .B1(n31), .Y(n30));
sg13g2_nor2_2 U21 (.A(n20), .B(n902), .Y(n31));
sg13g2_nand3_1 U22 (.A(n410), .B(n134), .C(n409), .Y(n779));
sg13g2_nand2_2 U23 (.A(data_i_85_), .B(n8), .Y(n607));
sg13g2_o21ai_1 U24 (.A1(n8), .A2(n344), .B1(n345), .Y(n754));
sg13g2_o21ai_1 U25 (.A1(n8), .A2(n256), .B1(n257), .Y(n730));
sg13g2_o21ai_1 U26 (.A1(n8), .A2(n36), .B1(n37), .Y(n670));
sg13g2_a21oi_2 U27 (.A1(outy_29_), .A2(n11), .B1(n38), .Y(n37));
sg13g2_nor2_2 U28 (.A(n14), .B(n310), .Y(n38));
sg13g2_o21ai_1 U29 (.A1(n15), .A2(n40), .B1(n41), .Y(n671));
sg13g2_a21oi_2 U30 (.A1(outy_29_), .A2(n18), .B1(n42), .Y(n41));
sg13g2_nor2_2 U31 (.A(n20), .B(n310), .Y(n42));
sg13g2_inv_4 U32 (.A(outx_25_), .Y(n39));
sg13g2_inv_4 U33 (.A(n39), .Y(n149));
sg13g2_a21oi_2 U34 (.A1(outx_28_), .A2(n4), .B1(n45), .Y(n44));
sg13g2_inv_4 U35 (.A(outy_13_), .Y(n211));
sg13g2_o21ai_1 U36 (.A1(n8), .A2(n47), .B1(n48), .Y(n673));
sg13g2_a21oi_2 U37 (.A1(outy_28_), .A2(n11), .B1(n49), .Y(n48));
sg13g2_nor2_2 U38 (.A(n14), .B(n50), .Y(n49));
sg13g2_o21ai_1 U39 (.A1(n15), .A2(n51), .B1(n52), .Y(n674));
sg13g2_a21oi_2 U40 (.A1(outy_28_), .A2(n18), .B1(n53), .Y(n52));
sg13g2_nor2_2 U41 (.A(n20), .B(n50), .Y(n53));
sg13g2_inv_4 U42 (.A(outx_28_), .Y(n50));
sg13g2_inv_4 U43 (.A(n211), .Y(n299));
sg13g2_a21oi_2 U44 (.A1(outx_27_), .A2(n4), .B1(n56), .Y(n55));
sg13g2_inv_4 U45 (.A(outy_22_), .Y(n112));
sg13g2_o21ai_1 U46 (.A1(n8), .A2(n58), .B1(n59), .Y(n676));
sg13g2_a21oi_2 U47 (.A1(outy_27_), .A2(n11), .B1(n60), .Y(n59));
sg13g2_nor2_2 U48 (.A(n14), .B(n61), .Y(n60));
sg13g2_o21ai_1 U49 (.A1(n15), .A2(n62), .B1(n63), .Y(n677));
sg13g2_a21oi_2 U50 (.A1(outy_27_), .A2(n18), .B1(n64), .Y(n63));
sg13g2_nor2_2 U51 (.A(n20), .B(n61), .Y(n64));
sg13g2_inv_4 U52 (.A(outx_27_), .Y(n61));
sg13g2_o21ai_1 U53 (.A1(n1), .A2(n65), .B1(n66), .Y(n678));
sg13g2_a21oi_2 U54 (.A1(outx_26_), .A2(n4), .B1(n67), .Y(n66));
sg13g2_nor2_2 U55 (.A(n6), .B(n68), .Y(n67));
sg13g2_o21ai_1 U56 (.A1(n8), .A2(n69), .B1(n70), .Y(n679));
sg13g2_a21oi_2 U57 (.A1(outy_26_), .A2(n11), .B1(n71), .Y(n70));
sg13g2_nor2_2 U58 (.A(n14), .B(n72), .Y(n71));
sg13g2_o21ai_1 U59 (.A1(n15), .A2(n73), .B1(n74), .Y(n680));
sg13g2_a21oi_2 U60 (.A1(outy_26_), .A2(n18), .B1(n75), .Y(n74));
sg13g2_nor2_2 U61 (.A(n20), .B(n72), .Y(n75));
sg13g2_inv_4 U62 (.A(outx_26_), .Y(n72));
sg13g2_o21ai_1 U63 (.A1(n1), .A2(n76), .B1(n77), .Y(n681));
sg13g2_a21oi_2 U64 (.A1(n149), .A2(n4), .B1(n78), .Y(n77));
sg13g2_nor2_2 U65 (.A(n6), .B(n79), .Y(n78));
sg13g2_nand2_2 U66 (.A(n662), .B(state_0_), .Y(n361));
sg13g2_a21oi_2 U67 (.A1(outy_25_), .A2(n11), .B1(n82), .Y(n81));
sg13g2_nor2_2 U68 (.A(n14), .B(n83), .Y(n82));
sg13g2_nand3_1 U69 (.A(n408), .B(n233), .C(n407), .Y(n778));
sg13g2_a21oi_2 U70 (.A1(outy_25_), .A2(n18), .B1(n86), .Y(n85));
sg13g2_nor2_2 U71 (.A(n20), .B(n83), .Y(n86));
sg13g2_inv_4 U72 (.A(outx_25_), .Y(n83));
sg13g2_o21ai_1 U73 (.A1(n1), .A2(n87), .B1(n88), .Y(n684));
sg13g2_a21oi_2 U74 (.A1(outx_24_), .A2(n4), .B1(n89), .Y(n88));
sg13g2_nand2_2 U75 (.A(n661), .B(state_1_), .Y(n355));
sg13g2_o21ai_1 U76 (.A1(n8), .A2(n91), .B1(n92), .Y(n685));
sg13g2_a21oi_2 U77 (.A1(outy_24_), .A2(n11), .B1(n93), .Y(n92));
sg13g2_nor2_2 U78 (.A(n14), .B(n94), .Y(n93));
sg13g2_o21ai_1 U79 (.A1(n15), .A2(n95), .B1(n96), .Y(n686));
sg13g2_a21oi_2 U80 (.A1(outy_24_), .A2(n18), .B1(n97), .Y(n96));
sg13g2_nor2_2 U81 (.A(n20), .B(n94), .Y(n97));
sg13g2_inv_4 U82 (.A(outx_24_), .Y(n94));
sg13g2_o21ai_1 U83 (.A1(n1), .A2(n98), .B1(n99), .Y(n687));
sg13g2_a21oi_2 U84 (.A1(outx_23_), .A2(n4), .B1(n100), .Y(n99));
sg13g2_nor2_2 U85 (.A(n6), .B(n101), .Y(n100));
sg13g2_o21ai_1 U86 (.A1(n8), .A2(n102), .B1(n103), .Y(n688));
sg13g2_a21oi_2 U87 (.A1(outy_23_), .A2(n11), .B1(n104), .Y(n103));
sg13g2_nor2_2 U88 (.A(n14), .B(n105), .Y(n104));
sg13g2_o21ai_1 U89 (.A1(n15), .A2(n106), .B1(n107), .Y(n689));
sg13g2_a21oi_2 U90 (.A1(outy_23_), .A2(n18), .B1(n108), .Y(n107));
sg13g2_nor2_2 U91 (.A(n20), .B(n105), .Y(n108));
sg13g2_inv_4 U92 (.A(outx_23_), .Y(n105));
sg13g2_nand3_1 U93 (.A(n426), .B(n908), .C(n425), .Y(n787));
sg13g2_a21oi_2 U94 (.A1(outx_22_), .A2(n4), .B1(n111), .Y(n110));
sg13g2_nor2_2 U95 (.A(n902), .B(n369), .Y(n903));
sg13g2_o21ai_1 U96 (.A1(n8), .A2(n113), .B1(n114), .Y(n691));
sg13g2_a21oi_2 U97 (.A1(n11), .A2(outy_22_), .B1(n115), .Y(n114));
sg13g2_nor2_2 U98 (.A(n14), .B(n116), .Y(n115));
sg13g2_o21ai_1 U99 (.A1(n15), .A2(n117), .B1(n118), .Y(n692));
sg13g2_a21oi_2 U100 (.A1(outy_22_), .A2(n18), .B1(n119), .Y(n118));
sg13g2_nor2_2 U101 (.A(n20), .B(n116), .Y(n119));
sg13g2_inv_4 U102 (.A(outx_22_), .Y(n116));
sg13g2_nand2_2 U103 (.A(n901), .B(n22), .Y(n666));
sg13g2_a21oi_2 U104 (.A1(outx_21_), .A2(n4), .B1(n122), .Y(n121));
sg13g2_nand4_1 U105 (.A(n637), .B(n638), .C(n639), .D(n640), .Y(mix_word_14_));
sg13g2_o21ai_1 U106 (.A1(n8), .A2(n124), .B1(n125), .Y(n694));
sg13g2_a21oi_2 U107 (.A1(n11), .A2(outy_21_), .B1(n126), .Y(n125));
sg13g2_nor2_2 U108 (.A(n14), .B(n127), .Y(n126));
sg13g2_o21ai_1 U109 (.A1(n15), .A2(n128), .B1(n129), .Y(n695));
sg13g2_a21oi_2 U110 (.A1(outy_21_), .A2(n18), .B1(n130), .Y(n129));
sg13g2_nor2_2 U111 (.A(n20), .B(n127), .Y(n130));
sg13g2_inv_4 U112 (.A(outx_21_), .Y(n127));
sg13g2_nand4_1 U113 (.A(n593), .B(n594), .C(n595), .D(n596), .Y(mix_word_24_));
sg13g2_a21oi_2 U114 (.A1(outx_20_), .A2(n4), .B1(n133), .Y(n132));
sg13g2_nor2_2 U115 (.A(n662), .B(n661), .Y(next_ready_o));
sg13g2_nor2_2 U116 (.A(n310), .B(n369), .Y(n889));
sg13g2_a21oi_2 U117 (.A1(outy_20_), .A2(n11), .B1(n137), .Y(n136));
sg13g2_nor2_2 U118 (.A(n14), .B(n138), .Y(n137));
sg13g2_nor2_2 U119 (.A(n889), .B(n34), .Y(n33));
sg13g2_a21oi_2 U120 (.A1(outy_20_), .A2(n18), .B1(n141), .Y(n140));
sg13g2_nor2_2 U121 (.A(n20), .B(n138), .Y(n141));
sg13g2_inv_4 U122 (.A(outx_20_), .Y(n138));
sg13g2_inv_4 U123 (.A(outx_29_), .Y(n310));
sg13g2_inv_4 U124 (.A(n4), .Y(n369));
sg13g2_nor2_2 U125 (.A(n6), .B(n893), .Y(n34));
sg13g2_nor2_2 U126 (.A(n905), .B(decrypt_i), .Y(n370));
sg13g2_a21oi_2 U127 (.A1(outy_19_), .A2(n11), .B1(n148), .Y(n147));
sg13g2_nor2_2 U128 (.A(n14), .B(n899), .Y(n148));
sg13g2_nor2_2 U129 (.A(n530), .B(n887), .Y(n433));
sg13g2_a21oi_2 U130 (.A1(outy_19_), .A2(n18), .B1(n152), .Y(n151));
sg13g2_nor2_2 U131 (.A(n20), .B(n899), .Y(n152));
sg13g2_inv_4 U132 (.A(outy_23_), .Y(n101));
sg13g2_inv_4 U133 (.A(outy_4_), .Y(n890));
sg13g2_a21oi_2 U134 (.A1(outx_18_), .A2(n4), .B1(n155), .Y(n154));
sg13g2_nor2_2 U135 (.A(n6), .B(n156), .Y(n155));
sg13g2_o21ai_1 U136 (.A1(n8), .A2(n157), .B1(n158), .Y(n703));
sg13g2_a21oi_2 U137 (.A1(outy_18_), .A2(n11), .B1(n159), .Y(n158));
sg13g2_nor2_2 U138 (.A(n14), .B(n160), .Y(n159));
sg13g2_o21ai_1 U139 (.A1(n15), .A2(n161), .B1(n162), .Y(n704));
sg13g2_a21oi_2 U140 (.A1(outy_18_), .A2(n18), .B1(n163), .Y(n162));
sg13g2_nor2_2 U141 (.A(n20), .B(n160), .Y(n163));
sg13g2_inv_4 U142 (.A(outx_18_), .Y(n160));
sg13g2_o21ai_1 U143 (.A1(n1), .A2(n164), .B1(n165), .Y(n705));
sg13g2_a21oi_2 U144 (.A1(outx_17_), .A2(n4), .B1(n166), .Y(n165));
sg13g2_nor2_2 U145 (.A(n6), .B(n167), .Y(n166));
sg13g2_nor2_2 U146 (.A(n123), .B(n6), .Y(n122));
sg13g2_a21oi_2 U147 (.A1(outy_17_), .A2(n11), .B1(n170), .Y(n169));
sg13g2_nor2_2 U148 (.A(n14), .B(n171), .Y(n170));
sg13g2_o21ai_1 U149 (.A1(n15), .A2(n172), .B1(n173), .Y(n707));
sg13g2_a21oi_2 U150 (.A1(outy_17_), .A2(n18), .B1(n174), .Y(n173));
sg13g2_nor2_2 U151 (.A(n20), .B(n171), .Y(n174));
sg13g2_inv_4 U152 (.A(outx_17_), .Y(n171));
sg13g2_inv_4 U153 (.A(outy_3_), .Y(n321));
sg13g2_a21oi_2 U154 (.A1(outx_16_), .A2(n4), .B1(n177), .Y(n176));
sg13g2_nor2_2 U155 (.A(n6), .B(n178), .Y(n177));
sg13g2_o21ai_1 U156 (.A1(n8), .A2(n179), .B1(n180), .Y(n709));
sg13g2_a21oi_2 U157 (.A1(outy_16_), .A2(n11), .B1(n181), .Y(n180));
sg13g2_nor2_2 U158 (.A(n14), .B(n182), .Y(n181));
sg13g2_o21ai_1 U159 (.A1(n15), .A2(n183), .B1(n184), .Y(n710));
sg13g2_a21oi_2 U160 (.A1(outy_16_), .A2(n18), .B1(n185), .Y(n184));
sg13g2_nor2_2 U161 (.A(n20), .B(n182), .Y(n185));
sg13g2_inv_4 U162 (.A(outx_16_), .Y(n182));
sg13g2_o21ai_1 U163 (.A1(n1), .A2(n186), .B1(n187), .Y(n711));
sg13g2_a21oi_2 U164 (.A1(outx_15_), .A2(n4), .B1(n188), .Y(n187));
sg13g2_nor2_2 U165 (.A(n365), .B(n360), .Y(n18));
sg13g2_o21ai_1 U166 (.A1(n8), .A2(n190), .B1(n191), .Y(n712));
sg13g2_a21oi_2 U167 (.A1(outy_15_), .A2(n11), .B1(n192), .Y(n191));
sg13g2_nor2_2 U168 (.A(n14), .B(n193), .Y(n192));
sg13g2_o21ai_1 U169 (.A1(n15), .A2(n194), .B1(n195), .Y(n713));
sg13g2_a21oi_2 U170 (.A1(outy_15_), .A2(n18), .B1(n196), .Y(n195));
sg13g2_nor2_2 U171 (.A(n20), .B(n193), .Y(n196));
sg13g2_inv_4 U172 (.A(outx_15_), .Y(n193));
sg13g2_o21ai_1 U173 (.A1(n1), .A2(n197), .B1(n198), .Y(n714));
sg13g2_a21oi_2 U174 (.A1(outx_14_), .A2(n4), .B1(n199), .Y(n198));
sg13g2_a21oi_2 U175 (.A1(n18), .A2(outy_31_), .B1(n19), .Y(n17));
sg13g2_o21ai_1 U176 (.A1(n8), .A2(n201), .B1(n202), .Y(n715));
sg13g2_a21oi_2 U177 (.A1(outy_14_), .A2(n11), .B1(n203), .Y(n202));
sg13g2_nor2_2 U178 (.A(n14), .B(n204), .Y(n203));
sg13g2_o21ai_1 U179 (.A1(n15), .A2(n205), .B1(n206), .Y(n716));
sg13g2_a21oi_2 U180 (.A1(outy_14_), .A2(n18), .B1(n207), .Y(n206));
sg13g2_nor2_2 U181 (.A(n20), .B(n204), .Y(n207));
sg13g2_inv_4 U182 (.A(outx_14_), .Y(n204));
sg13g2_o21ai_1 U183 (.A1(n1), .A2(n142), .B1(n143), .Y(n699));
sg13g2_a21oi_2 U184 (.A1(outx_13_), .A2(n4), .B1(n210), .Y(n209));
sg13g2_nor2_2 U185 (.A(n6), .B(n891), .Y(n210));
sg13g2_o21ai_1 U186 (.A1(n8), .A2(n212), .B1(n213), .Y(n718));
sg13g2_a21oi_2 U187 (.A1(n11), .A2(n299), .B1(n214), .Y(n213));
sg13g2_nor2_2 U188 (.A(n14), .B(n215), .Y(n214));
sg13g2_o21ai_1 U189 (.A1(n15), .A2(n216), .B1(n217), .Y(n719));
sg13g2_a21oi_2 U190 (.A1(n18), .A2(n299), .B1(n218), .Y(n217));
sg13g2_nor2_2 U191 (.A(n20), .B(n215), .Y(n218));
sg13g2_inv_4 U192 (.A(outx_13_), .Y(n215));
sg13g2_o21ai_1 U193 (.A1(n15), .A2(n150), .B1(n151), .Y(n701));
sg13g2_a21oi_2 U194 (.A1(outx_12_), .A2(n4), .B1(n221), .Y(n220));
sg13g2_nand3_1 U195 (.A(n424), .B(n909), .C(n423), .Y(n786));
sg13g2_inv_4 U196 (.A(outy_21_), .Y(n123));
sg13g2_a21oi_2 U197 (.A1(outy_12_), .A2(n11), .B1(n225), .Y(n224));
sg13g2_nor2_2 U198 (.A(n14), .B(n226), .Y(n225));
sg13g2_o21ai_1 U199 (.A1(n15), .A2(n227), .B1(n228), .Y(n722));
sg13g2_a21oi_2 U200 (.A1(outy_12_), .A2(n18), .B1(n229), .Y(n228));
sg13g2_inv_4 U201 (.A(outy_13_), .Y(n891));
sg13g2_inv_4 U202 (.A(outx_12_), .Y(n226));
sg13g2_nor2_2 U203 (.A(n6), .B(n200), .Y(n199));
sg13g2_a21oi_2 U204 (.A1(outx_11_), .A2(n4), .B1(n232), .Y(n231));
sg13g2_o21ai_1 U205 (.A1(n8), .A2(n146), .B1(n147), .Y(n700));
sg13g2_o21ai_1 U206 (.A1(n8), .A2(n234), .B1(n235), .Y(n724));
sg13g2_a21oi_2 U207 (.A1(n11), .A2(outy_11_), .B1(n236), .Y(n235));
sg13g2_nor2_2 U208 (.A(n14), .B(n237), .Y(n236));
sg13g2_o21ai_1 U209 (.A1(n15), .A2(n238), .B1(n239), .Y(n725));
sg13g2_a21oi_2 U210 (.A1(n18), .A2(outy_11_), .B1(n240), .Y(n239));
sg13g2_nor2_2 U211 (.A(n20), .B(n237), .Y(n240));
sg13g2_inv_4 U212 (.A(outx_11_), .Y(n237));
sg13g2_o21ai_1 U213 (.A1(n1), .A2(n241), .B1(n242), .Y(n726));
sg13g2_a21oi_2 U214 (.A1(outx_10_), .A2(n4), .B1(n243), .Y(n242));
sg13g2_nor2_2 U215 (.A(n6), .B(n244), .Y(n243));
sg13g2_o21ai_1 U216 (.A1(n8), .A2(n245), .B1(n246), .Y(n727));
sg13g2_a21oi_2 U217 (.A1(outy_10_), .A2(n11), .B1(n247), .Y(n246));
sg13g2_nor2_2 U218 (.A(n14), .B(n248), .Y(n247));
sg13g2_o21ai_1 U219 (.A1(n15), .A2(n249), .B1(n250), .Y(n728));
sg13g2_a21oi_2 U220 (.A1(outy_10_), .A2(n18), .B1(n251), .Y(n250));
sg13g2_nor2_2 U221 (.A(n20), .B(n248), .Y(n251));
sg13g2_inv_4 U222 (.A(outx_10_), .Y(n248));
sg13g2_o21ai_1 U223 (.A1(n1), .A2(n252), .B1(n253), .Y(n729));
sg13g2_a21oi_2 U224 (.A1(outx_9_), .A2(n4), .B1(n254), .Y(n253));
sg13g2_nor2_2 U225 (.A(n6), .B(n255), .Y(n254));
sg13g2_o21ai_1 U226 (.A1(n1), .A2(n285), .B1(n286), .Y(n738));
sg13g2_a21oi_2 U227 (.A1(outy_9_), .A2(n11), .B1(n258), .Y(n257));
sg13g2_nand3_1 U228 (.A(n412), .B(n910), .C(n411), .Y(n780));
sg13g2_nand3_1 U229 (.A(n428), .B(n911), .C(n427), .Y(n788));
sg13g2_a21oi_2 U230 (.A1(outy_9_), .A2(n18), .B1(n262), .Y(n261));
sg13g2_nor2_2 U231 (.A(n20), .B(n259), .Y(n262));
sg13g2_inv_4 U232 (.A(outx_9_), .Y(n259));
sg13g2_o21ai_1 U233 (.A1(n15), .A2(n260), .B1(n261), .Y(n731));
sg13g2_a21oi_2 U234 (.A1(outx_8_), .A2(n4), .B1(n265), .Y(n264));
sg13g2_nor2_2 U235 (.A(n6), .B(n266), .Y(n265));
sg13g2_o21ai_1 U236 (.A1(n8), .A2(n267), .B1(n268), .Y(n733));
sg13g2_a21oi_2 U237 (.A1(outy_8_), .A2(n11), .B1(n269), .Y(n268));
sg13g2_nor2_2 U238 (.A(n14), .B(n270), .Y(n269));
sg13g2_o21ai_1 U239 (.A1(n15), .A2(n271), .B1(n272), .Y(n734));
sg13g2_a21oi_2 U240 (.A1(outy_8_), .A2(n18), .B1(n273), .Y(n272));
sg13g2_nor2_2 U241 (.A(n20), .B(n270), .Y(n273));
sg13g2_inv_4 U242 (.A(outx_8_), .Y(n270));
sg13g2_o21ai_1 U243 (.A1(n1), .A2(n274), .B1(n275), .Y(n735));
sg13g2_a21oi_2 U244 (.A1(outx_7_), .A2(n4), .B1(n276), .Y(n275));
sg13g2_nor2_2 U245 (.A(n6), .B(n277), .Y(n276));
sg13g2_o21ai_1 U246 (.A1(n8), .A2(n278), .B1(n279), .Y(n736));
sg13g2_a21oi_2 U247 (.A1(outy_7_), .A2(n11), .B1(n280), .Y(n279));
sg13g2_nor2_2 U248 (.A(n14), .B(n281), .Y(n280));
sg13g2_o21ai_1 U249 (.A1(n15), .A2(n282), .B1(n283), .Y(n737));
sg13g2_a21oi_2 U250 (.A1(outy_7_), .A2(n18), .B1(n284), .Y(n283));
sg13g2_nor2_2 U251 (.A(n20), .B(n281), .Y(n284));
sg13g2_inv_4 U252 (.A(outx_7_), .Y(n281));
sg13g2_nor2_2 U253 (.A(n6), .B(n145), .Y(n144));
sg13g2_a21oi_2 U254 (.A1(outx_6_), .A2(n4), .B1(n287), .Y(n286));
sg13g2_nor2_2 U255 (.A(n900), .B(n144), .Y(n143));
sg13g2_o21ai_1 U256 (.A1(n8), .A2(n289), .B1(n290), .Y(n739));
sg13g2_a21oi_2 U257 (.A1(outy_6_), .A2(n11), .B1(n291), .Y(n290));
sg13g2_nor2_2 U258 (.A(n14), .B(n292), .Y(n291));
sg13g2_o21ai_1 U259 (.A1(n15), .A2(n293), .B1(n294), .Y(n740));
sg13g2_a21oi_2 U260 (.A1(outy_6_), .A2(n18), .B1(n295), .Y(n294));
sg13g2_nor2_2 U261 (.A(n20), .B(n292), .Y(n295));
sg13g2_inv_4 U262 (.A(outx_6_), .Y(n292));
sg13g2_nand3_1 U263 (.A(n432), .B(n912), .C(n431), .Y(n790));
sg13g2_a21oi_2 U264 (.A1(outx_5_), .A2(n4), .B1(n298), .Y(n297));
sg13g2_inv_4 U265 (.A(outy_19_), .Y(n145));
sg13g2_o21ai_1 U266 (.A1(n8), .A2(n300), .B1(n301), .Y(n742));
sg13g2_a21oi_2 U267 (.A1(n11), .A2(n35), .B1(n302), .Y(n301));
sg13g2_nor2_2 U268 (.A(n14), .B(n303), .Y(n302));
sg13g2_o21ai_1 U269 (.A1(n15), .A2(n304), .B1(n305), .Y(n743));
sg13g2_a21oi_2 U270 (.A1(n35), .A2(n18), .B1(n306), .Y(n305));
sg13g2_nor2_2 U271 (.A(n20), .B(n303), .Y(n306));
sg13g2_inv_4 U272 (.A(outx_5_), .Y(n303));
sg13g2_inv_4 U273 (.A(outy_5_), .Y(n892));
sg13g2_a21oi_2 U274 (.A1(outx_4_), .A2(n4), .B1(n309), .Y(n308));
sg13g2_nor2_2 U275 (.A(n903), .B(n23), .Y(n22));
sg13g2_o21ai_1 U276 (.A1(n8), .A2(n168), .B1(n169), .Y(n706));
sg13g2_a21oi_2 U277 (.A1(outy_4_), .A2(n11), .B1(n313), .Y(n312));
sg13g2_nor2_2 U278 (.A(n14), .B(n314), .Y(n313));
sg13g2_nor2_2 U279 (.A(n6), .B(n7), .Y(n5));
sg13g2_a21oi_2 U280 (.A1(outy_4_), .A2(n18), .B1(n317), .Y(n316));
sg13g2_nor2_2 U281 (.A(n20), .B(n314), .Y(n317));
sg13g2_inv_4 U282 (.A(outx_4_), .Y(n314));
sg13g2_inv_4 U283 (.A(outy_31_), .Y(n7));
sg13g2_a21oi_2 U284 (.A1(outx_3_), .A2(n4), .B1(n320), .Y(n319));
sg13g2_inv_4 U285 (.A(outy_29_), .Y(n893));
sg13g2_o21ai_1 U286 (.A1(n8), .A2(n322), .B1(n323), .Y(n748));
sg13g2_a21oi_2 U287 (.A1(n11), .A2(outy_3_), .B1(n324), .Y(n323));
sg13g2_nor2_2 U288 (.A(n14), .B(n325), .Y(n324));
sg13g2_o21ai_1 U289 (.A1(n15), .A2(n326), .B1(n327), .Y(n749));
sg13g2_a21oi_2 U290 (.A1(outy_3_), .A2(n18), .B1(n328), .Y(n327));
sg13g2_nor2_2 U291 (.A(n20), .B(n325), .Y(n328));
sg13g2_inv_4 U292 (.A(outx_3_), .Y(n325));
sg13g2_o21ai_1 U293 (.A1(n1), .A2(n329), .B1(n330), .Y(n750));
sg13g2_a21oi_2 U294 (.A1(outx_2_), .A2(n4), .B1(n331), .Y(n330));
sg13g2_nor2_2 U295 (.A(n6), .B(n332), .Y(n331));
sg13g2_o21ai_1 U296 (.A1(n8), .A2(n333), .B1(n334), .Y(n751));
sg13g2_a21oi_2 U297 (.A1(outy_2_), .A2(n11), .B1(n335), .Y(n334));
sg13g2_nor2_2 U298 (.A(n14), .B(n336), .Y(n335));
sg13g2_o21ai_1 U299 (.A1(n15), .A2(n337), .B1(n338), .Y(n752));
sg13g2_a21oi_2 U300 (.A1(outy_2_), .A2(n18), .B1(n339), .Y(n338));
sg13g2_nor2_2 U301 (.A(n20), .B(n336), .Y(n339));
sg13g2_inv_4 U302 (.A(outx_2_), .Y(n336));
sg13g2_o21ai_1 U303 (.A1(n1), .A2(n340), .B1(n341), .Y(n753));
sg13g2_a21oi_2 U304 (.A1(outx_1_), .A2(n4), .B1(n342), .Y(n341));
sg13g2_nor2_2 U305 (.A(n6), .B(n343), .Y(n342));
sg13g2_nand2_2 U306 (.A(data_i_71_), .B(n8), .Y(n543));
sg13g2_a21oi_2 U307 (.A1(outy_1_), .A2(n11), .B1(n346), .Y(n345));
sg13g2_nor2_2 U308 (.A(n14), .B(n347), .Y(n346));
sg13g2_o21ai_1 U309 (.A1(n15), .A2(n348), .B1(n349), .Y(n755));
sg13g2_a21oi_2 U310 (.A1(outy_1_), .A2(n18), .B1(n350), .Y(n349));
sg13g2_nor2_2 U311 (.A(n20), .B(n347), .Y(n350));
sg13g2_inv_4 U312 (.A(outx_1_), .Y(n347));
sg13g2_nor2_2 U313 (.A(n14), .B(n259), .Y(n258));
sg13g2_a21oi_2 U314 (.A1(outx_0_), .A2(n4), .B1(n353), .Y(n352));
sg13g2_nor2_2 U315 (.A(n6), .B(n354), .Y(n353));
sg13g2_nand2_2 U316 (.A(decrypt_i), .B(n1), .Y(n6));
sg13g2_nor2_2 U317 (.A(n355), .B(decrypt_i), .Y(n4));
sg13g2_o21ai_1 U318 (.A1(n8), .A2(n356), .B1(n357), .Y(n757));
sg13g2_a21oi_2 U319 (.A1(outy_0_), .A2(n11), .B1(n358), .Y(n357));
sg13g2_nor2_2 U320 (.A(n14), .B(n359), .Y(n358));
sg13g2_nand2_2 U321 (.A(n8), .B(n360), .Y(n14));
sg13g2_nor2_2 U322 (.A(n361), .B(n360), .Y(n11));
sg13g2_o21ai_1 U323 (.A1(n15), .A2(n362), .B1(n363), .Y(n758));
sg13g2_a21oi_2 U324 (.A1(outy_0_), .A2(n18), .B1(n364), .Y(n363));
sg13g2_nor2_2 U325 (.A(n20), .B(n359), .Y(n364));
sg13g2_inv_4 U326 (.A(outx_0_), .Y(n359));
sg13g2_nand2_2 U327 (.A(n15), .B(n360), .Y(n20));
sg13g2_o21ai_1 U328 (.A1(n1), .A2(n296), .B1(n297), .Y(n741));
sg13g2_inv_4 U329 (.A(decrypt_i), .Y(n360));
sg13g2_nand3_1 U330 (.A(n422), .B(n913), .C(n421), .Y(n785));
sg13g2_nand2_2 U331 (.A(data_o_0_), .B(n906), .Y(n368));
sg13g2_nand2_2 U332 (.A(n370), .B(outx_0_), .Y(n367));
sg13g2_inv_4 U333 (.A(outy_0_), .Y(n354));
sg13g2_nand3_1 U334 (.A(n420), .B(n914), .C(n419), .Y(n784));
sg13g2_nand2_2 U335 (.A(data_o_1_), .B(n907), .Y(n372));
sg13g2_nand2_2 U336 (.A(n370), .B(outx_1_), .Y(n371));
sg13g2_inv_4 U337 (.A(outy_1_), .Y(n343));
sg13g2_nand3_1 U338 (.A(n418), .B(n915), .C(n417), .Y(n783));
sg13g2_nand2_2 U339 (.A(data_o_2_), .B(n904), .Y(n374));
sg13g2_nand2_2 U340 (.A(n370), .B(outx_2_), .Y(n373));
sg13g2_inv_4 U341 (.A(outy_2_), .Y(n332));
sg13g2_nand3_1 U342 (.A(n416), .B(n916), .C(n415), .Y(n782));
sg13g2_nand2_2 U343 (.A(data_o_3_), .B(n907), .Y(n376));
sg13g2_nand2_2 U344 (.A(n370), .B(outx_3_), .Y(n375));
sg13g2_nor2_2 U345 (.A(n6), .B(n189), .Y(n188));
sg13g2_nand3_1 U346 (.A(n414), .B(n917), .C(n413), .Y(n781));
sg13g2_nand2_2 U347 (.A(data_o_4_), .B(n907), .Y(n378));
sg13g2_nand2_2 U348 (.A(n370), .B(outx_4_), .Y(n377));
sg13g2_inv_4 U349 (.A(outy_15_), .Y(n189));
sg13g2_nand3_1 U350 (.A(n406), .B(n918), .C(n405), .Y(n777));
sg13g2_nand2_2 U351 (.A(data_o_5_), .B(n906), .Y(n380));
sg13g2_nand2_2 U352 (.A(n370), .B(outx_5_), .Y(n379));
sg13g2_nand2_2 U353 (.A(data_i_63_), .B(n1), .Y(n564));
sg13g2_nand3_1 U354 (.A(n404), .B(n919), .C(n403), .Y(n776));
sg13g2_nand2_2 U355 (.A(data_o_6_), .B(n906), .Y(n382));
sg13g2_nand2_2 U356 (.A(n370), .B(outx_6_), .Y(n381));
sg13g2_inv_4 U357 (.A(outy_6_), .Y(n288));
sg13g2_nand3_1 U358 (.A(n402), .B(n920), .C(n401), .Y(n775));
sg13g2_nand2_2 U359 (.A(data_o_7_), .B(n905), .Y(n384));
sg13g2_nand2_2 U360 (.A(n370), .B(outx_7_), .Y(n383));
sg13g2_inv_4 U361 (.A(outy_7_), .Y(n277));
sg13g2_nand3_1 U362 (.A(n400), .B(n921), .C(n399), .Y(n774));
sg13g2_nand2_2 U363 (.A(data_o_8_), .B(n905), .Y(n386));
sg13g2_nand2_2 U364 (.A(n370), .B(outx_8_), .Y(n385));
sg13g2_inv_4 U365 (.A(outy_8_), .Y(n266));
sg13g2_nand3_1 U366 (.A(n398), .B(n922), .C(n397), .Y(n773));
sg13g2_nand2_2 U367 (.A(data_o_9_), .B(n906), .Y(n388));
sg13g2_nand2_2 U368 (.A(n370), .B(outx_9_), .Y(n387));
sg13g2_inv_4 U369 (.A(outy_9_), .Y(n255));
sg13g2_nand3_1 U370 (.A(n396), .B(n923), .C(n395), .Y(n772));
sg13g2_nand2_2 U371 (.A(data_o_10_), .B(n907), .Y(n390));
sg13g2_nand2_2 U372 (.A(n370), .B(outx_10_), .Y(n389));
sg13g2_inv_4 U373 (.A(outy_10_), .Y(n244));
sg13g2_nand2_2 U374 (.A(data_i_93_), .B(n8), .Y(n575));
sg13g2_nand2_2 U375 (.A(data_o_11_), .B(n905), .Y(n392));
sg13g2_nand2_2 U376 (.A(n370), .B(outx_11_), .Y(n391));
sg13g2_nand3_1 U377 (.A(n394), .B(n924), .C(n393), .Y(n771));
sg13g2_nand3_1 U378 (.A(n390), .B(n925), .C(n389), .Y(n769));
sg13g2_nand2_2 U379 (.A(data_o_12_), .B(n904), .Y(n394));
sg13g2_nand2_2 U380 (.A(n370), .B(outx_12_), .Y(n393));
sg13g2_inv_4 U381 (.A(outy_12_), .Y(n222));
sg13g2_nand3_1 U382 (.A(n388), .B(n926), .C(n387), .Y(n768));
sg13g2_nand2_2 U383 (.A(data_o_13_), .B(n907), .Y(n396));
sg13g2_nand2_2 U384 (.A(n370), .B(outx_13_), .Y(n395));
sg13g2_nand3_1 U385 (.A(n386), .B(n927), .C(n385), .Y(n767));
sg13g2_nand3_1 U386 (.A(n384), .B(n928), .C(n383), .Y(n766));
sg13g2_nand2_2 U387 (.A(data_o_14_), .B(n905), .Y(n398));
sg13g2_nand2_2 U388 (.A(n370), .B(outx_14_), .Y(n397));
sg13g2_inv_4 U389 (.A(outy_14_), .Y(n200));
sg13g2_nand3_1 U390 (.A(n382), .B(n929), .C(n381), .Y(n765));
sg13g2_nand2_2 U391 (.A(data_o_15_), .B(n906), .Y(n400));
sg13g2_nand2_2 U392 (.A(n370), .B(outx_15_), .Y(n399));
sg13g2_nand2_2 U393 (.A(data_i_39_), .B(n1), .Y(n544));
sg13g2_nand3_1 U394 (.A(n380), .B(n930), .C(n379), .Y(n764));
sg13g2_nand2_2 U395 (.A(data_o_16_), .B(n905), .Y(n402));
sg13g2_nand2_2 U396 (.A(n370), .B(outx_16_), .Y(n401));
sg13g2_inv_4 U397 (.A(outy_16_), .Y(n178));
sg13g2_nand3_1 U398 (.A(n378), .B(n931), .C(n377), .Y(n763));
sg13g2_nand2_2 U399 (.A(data_o_17_), .B(n905), .Y(n404));
sg13g2_nand2_2 U400 (.A(n370), .B(outx_17_), .Y(n403));
sg13g2_inv_4 U401 (.A(outy_17_), .Y(n167));
sg13g2_nand3_1 U402 (.A(n376), .B(n932), .C(n375), .Y(n762));
sg13g2_nand2_2 U403 (.A(data_o_18_), .B(n907), .Y(n406));
sg13g2_nand2_2 U404 (.A(n370), .B(outx_18_), .Y(n405));
sg13g2_inv_4 U405 (.A(outy_18_), .Y(n156));
sg13g2_nand2_2 U406 (.A(data_i_13_), .B(next_ready_o), .Y(n641));
sg13g2_nand2_2 U407 (.A(data_o_19_), .B(n905), .Y(n408));
sg13g2_nand2_2 U408 (.A(n370), .B(outx_19_), .Y(n407));
sg13g2_nand3_1 U409 (.A(n374), .B(n933), .C(n373), .Y(n761));
sg13g2_nand2_2 U410 (.A(data_i_21_), .B(next_ready_o), .Y(n605));
sg13g2_nand2_2 U411 (.A(data_o_20_), .B(n905), .Y(n410));
sg13g2_nand2_2 U412 (.A(n370), .B(outx_20_), .Y(n409));
sg13g2_nand3_1 U413 (.A(n372), .B(n934), .C(n371), .Y(n760));
sg13g2_nand2_2 U414 (.A(data_i_117_), .B(n15), .Y(n606));
sg13g2_nand2_2 U415 (.A(data_o_21_), .B(n907), .Y(n412));
sg13g2_nand2_2 U416 (.A(n370), .B(outx_21_), .Y(n411));
sg13g2_nand3_1 U417 (.A(n368), .B(n935), .C(n367), .Y(n759));
sg13g2_inv_1 U418 (.A(n366), .Y(n936));
sg13g2_nand2_2 U419 (.A(data_o_22_), .B(n905), .Y(n414));
sg13g2_nand2_2 U420 (.A(n370), .B(outx_22_), .Y(n413));
sg13g2_o21ai_1 U421 (.A1(n1), .A2(n230), .B1(n231), .Y(n723));
sg13g2_nand2_1 U422 (.A(outy_31_), .B(n936), .Y(n912));
sg13g2_nand2_2 U423 (.A(data_o_23_), .B(n904), .Y(n416));
sg13g2_nand2_2 U424 (.A(n370), .B(outx_23_), .Y(n415));
sg13g2_nand2_2 U425 (.A(data_i_109_), .B(n15), .Y(n642));
sg13g2_nand2_1 U426 (.A(outy_30_), .B(n936), .Y(n46));
sg13g2_nand2_2 U427 (.A(data_o_24_), .B(n905), .Y(n418));
sg13g2_nand2_2 U428 (.A(n370), .B(outx_24_), .Y(n417));
sg13g2_inv_4 U429 (.A(outy_24_), .Y(n90));
sg13g2_nand2_1 U430 (.A(outy_29_), .B(n936), .Y(n911));
sg13g2_nand2_2 U431 (.A(data_o_25_), .B(n904), .Y(n420));
sg13g2_nand2_2 U432 (.A(n370), .B(n149), .Y(n419));
sg13g2_inv_4 U433 (.A(outy_25_), .Y(n79));
sg13g2_nand2_1 U434 (.A(outy_28_), .B(n936), .Y(n908));
sg13g2_nand2_2 U435 (.A(data_o_26_), .B(n905), .Y(n422));
sg13g2_nand2_2 U436 (.A(n370), .B(outx_26_), .Y(n421));
sg13g2_inv_4 U437 (.A(outy_26_), .Y(n68));
sg13g2_nor2_2 U438 (.A(n222), .B(n6), .Y(n221));
sg13g2_nand2_2 U439 (.A(data_o_27_), .B(n907), .Y(n424));
sg13g2_nand2_2 U440 (.A(n370), .B(outx_27_), .Y(n423));
sg13g2_nand2_1 U441 (.A(outy_27_), .B(n936), .Y(n909));
sg13g2_nand2_2 U442 (.A(outy_28_), .B(n896), .Y(n894));
sg13g2_nand2_2 U443 (.A(data_o_28_), .B(n906), .Y(n426));
sg13g2_nand2_2 U444 (.A(n370), .B(outx_28_), .Y(n425));
sg13g2_nand2_1 U445 (.A(outy_26_), .B(n936), .Y(n913));
sg13g2_inv_4 U446 (.A(n894), .Y(n45));
sg13g2_nand2_2 U447 (.A(data_o_29_), .B(n907), .Y(n428));
sg13g2_nand2_2 U448 (.A(n370), .B(outx_29_), .Y(n427));
sg13g2_nand4_1 U449 (.A(n575), .B(n573), .C(n574), .D(n576), .Y(mix_word_29_));
sg13g2_nand3_1 U450 (.A(decrypt_i), .B(outy_27_), .C(n1), .Y(n895));
sg13g2_nand2_2 U451 (.A(data_o_30_), .B(n905), .Y(n430));
sg13g2_nand2_2 U452 (.A(n370), .B(outx_30_), .Y(n429));
sg13g2_inv_4 U453 (.A(outy_30_), .Y(n24));
sg13g2_nand2_1 U454 (.A(outy_25_), .B(n936), .Y(n914));
sg13g2_nand2_2 U455 (.A(data_o_31_), .B(n907), .Y(n432));
sg13g2_nand2_2 U456 (.A(n370), .B(outx_31_), .Y(n431));
sg13g2_inv_4 U457 (.A(n895), .Y(n56));
sg13g2_nand2_2 U458 (.A(n433), .B(decrypt_i), .Y(n366));
sg13g2_nand2_2 U459 (.A(outy_11_), .B(n896), .Y(n897));
sg13g2_o21ai_1 U460 (.A1(n351), .A2(n906), .B1(n434), .Y(n791));
sg13g2_nand2_2 U461 (.A(data_o_32_), .B(n907), .Y(n434));
sg13g2_nand2_1 U462 (.A(outy_24_), .B(n936), .Y(n915));
sg13g2_o21ai_1 U463 (.A1(n340), .A2(n906), .B1(n435), .Y(n792));
sg13g2_nand2_2 U464 (.A(data_o_33_), .B(n906), .Y(n435));
sg13g2_nand2_1 U465 (.A(outy_23_), .B(n936), .Y(n916));
sg13g2_o21ai_1 U466 (.A1(n329), .A2(n907), .B1(n436), .Y(n793));
sg13g2_nand2_2 U467 (.A(data_o_34_), .B(n906), .Y(n436));
sg13g2_nand2_1 U468 (.A(outy_22_), .B(n936), .Y(n917));
sg13g2_o21ai_1 U469 (.A1(n318), .A2(n906), .B1(n437), .Y(n794));
sg13g2_nand2_2 U470 (.A(data_o_35_), .B(n904), .Y(n437));
sg13g2_nand2_1 U471 (.A(outy_21_), .B(n936), .Y(n910));
sg13g2_o21ai_1 U472 (.A1(n307), .A2(n906), .B1(n438), .Y(n795));
sg13g2_nand2_2 U473 (.A(data_o_36_), .B(n904), .Y(n438));
sg13g2_nand2_1 U474 (.A(outy_20_), .B(n936), .Y(n134));
sg13g2_o21ai_1 U475 (.A1(n296), .A2(n907), .B1(n439), .Y(n796));
sg13g2_nand2_2 U476 (.A(data_o_37_), .B(n906), .Y(n439));
sg13g2_nand2_1 U477 (.A(outy_19_), .B(n936), .Y(n233));
sg13g2_o21ai_1 U478 (.A1(n285), .A2(n907), .B1(n440), .Y(n797));
sg13g2_nand2_2 U479 (.A(data_o_38_), .B(n904), .Y(n440));
sg13g2_nand2_1 U480 (.A(outy_18_), .B(n936), .Y(n918));
sg13g2_o21ai_1 U481 (.A1(n274), .A2(n907), .B1(n441), .Y(n798));
sg13g2_nand2_2 U482 (.A(data_o_39_), .B(n904), .Y(n441));
sg13g2_nand2_1 U483 (.A(outy_17_), .B(n936), .Y(n919));
sg13g2_o21ai_1 U484 (.A1(n263), .A2(n907), .B1(n442), .Y(n799));
sg13g2_nand2_2 U485 (.A(data_o_40_), .B(n907), .Y(n442));
sg13g2_nand2_1 U486 (.A(outy_16_), .B(n936), .Y(n920));
sg13g2_o21ai_1 U487 (.A1(n252), .A2(n907), .B1(n443), .Y(n800));
sg13g2_nand2_2 U488 (.A(data_o_41_), .B(n906), .Y(n443));
sg13g2_nand2_1 U489 (.A(outy_15_), .B(n936), .Y(n921));
sg13g2_o21ai_1 U490 (.A1(n241), .A2(n906), .B1(n444), .Y(n801));
sg13g2_nand2_2 U491 (.A(data_o_42_), .B(n904), .Y(n444));
sg13g2_nand2_1 U492 (.A(outy_14_), .B(n936), .Y(n922));
sg13g2_o21ai_1 U493 (.A1(n230), .A2(n906), .B1(n445), .Y(n802));
sg13g2_nand2_2 U494 (.A(data_o_43_), .B(n904), .Y(n445));
sg13g2_nand2_1 U495 (.A(n299), .B(n936), .Y(n923));
sg13g2_o21ai_1 U496 (.A1(n219), .A2(n904), .B1(n446), .Y(n803));
sg13g2_nand2_2 U497 (.A(data_o_44_), .B(n904), .Y(n446));
sg13g2_nand2_1 U498 (.A(outy_12_), .B(n936), .Y(n924));
sg13g2_o21ai_1 U499 (.A1(n208), .A2(n907), .B1(n447), .Y(n804));
sg13g2_nand2_2 U500 (.A(data_o_45_), .B(n905), .Y(n447));
sg13g2_nand2_1 U501 (.A(outy_11_), .B(n936), .Y(n57));
sg13g2_o21ai_1 U502 (.A1(n197), .A2(n906), .B1(n448), .Y(n805));
sg13g2_nand2_2 U503 (.A(data_o_46_), .B(n906), .Y(n448));
sg13g2_nand2_1 U504 (.A(outy_10_), .B(n936), .Y(n925));
sg13g2_o21ai_1 U505 (.A1(n186), .A2(n905), .B1(n449), .Y(n806));
sg13g2_nand2_2 U506 (.A(data_o_47_), .B(n907), .Y(n449));
sg13g2_nand2_1 U507 (.A(outy_9_), .B(n936), .Y(n926));
sg13g2_o21ai_1 U508 (.A1(n175), .A2(n904), .B1(n450), .Y(n807));
sg13g2_nand2_2 U509 (.A(data_o_48_), .B(n904), .Y(n450));
sg13g2_nand2_1 U510 (.A(outy_8_), .B(n936), .Y(n927));
sg13g2_o21ai_1 U511 (.A1(n164), .A2(n904), .B1(n451), .Y(n808));
sg13g2_nand2_2 U512 (.A(data_o_49_), .B(n906), .Y(n451));
sg13g2_nand2_1 U513 (.A(outy_7_), .B(n936), .Y(n928));
sg13g2_o21ai_1 U514 (.A1(n153), .A2(n906), .B1(n452), .Y(n809));
sg13g2_nand2_2 U515 (.A(data_o_50_), .B(n905), .Y(n452));
sg13g2_nand2_1 U516 (.A(outy_6_), .B(n936), .Y(n929));
sg13g2_o21ai_1 U517 (.A1(n142), .A2(n905), .B1(n453), .Y(n810));
sg13g2_nand2_2 U518 (.A(data_o_51_), .B(n906), .Y(n453));
sg13g2_nand2_1 U519 (.A(n35), .B(n936), .Y(n930));
sg13g2_o21ai_1 U520 (.A1(n131), .A2(n906), .B1(n454), .Y(n811));
sg13g2_nand2_2 U521 (.A(data_o_52_), .B(n907), .Y(n454));
sg13g2_nand2_1 U522 (.A(outy_4_), .B(n936), .Y(n931));
sg13g2_o21ai_1 U523 (.A1(n120), .A2(n907), .B1(n455), .Y(n812));
sg13g2_nand2_2 U524 (.A(data_o_53_), .B(n904), .Y(n455));
sg13g2_nand2_1 U525 (.A(outy_3_), .B(n936), .Y(n932));
sg13g2_o21ai_1 U526 (.A1(n109), .A2(n906), .B1(n456), .Y(n813));
sg13g2_nand2_2 U527 (.A(data_o_54_), .B(n904), .Y(n456));
sg13g2_nand2_1 U528 (.A(outy_2_), .B(n936), .Y(n933));
sg13g2_o21ai_1 U529 (.A1(n98), .A2(n905), .B1(n457), .Y(n814));
sg13g2_nand2_2 U530 (.A(data_o_55_), .B(n907), .Y(n457));
sg13g2_nand2_1 U531 (.A(outy_1_), .B(n936), .Y(n934));
sg13g2_o21ai_1 U532 (.A1(n87), .A2(n907), .B1(n458), .Y(n815));
sg13g2_nand2_2 U533 (.A(data_o_56_), .B(n906), .Y(n458));
sg13g2_nand2_1 U534 (.A(outy_0_), .B(n936), .Y(n935));
sg13g2_o21ai_1 U535 (.A1(n76), .A2(n905), .B1(n459), .Y(n816));
sg13g2_nand2_2 U536 (.A(data_o_57_), .B(n907), .Y(n459));
sg13g2_o21ai_1 U538 (.A1(n65), .A2(n904), .B1(n460), .Y(n817));
sg13g2_nand2_2 U539 (.A(data_o_58_), .B(n906), .Y(n460));
sg13g2_o21ai_1 U541 (.A1(n54), .A2(n906), .B1(n461), .Y(n818));
sg13g2_nand2_2 U542 (.A(data_o_59_), .B(n906), .Y(n461));
sg13g2_o21ai_1 U544 (.A1(n43), .A2(n906), .B1(n462), .Y(n819));
sg13g2_nand2_2 U545 (.A(data_o_60_), .B(n905), .Y(n462));
sg13g2_o21ai_1 U547 (.A1(n32), .A2(n907), .B1(n463), .Y(n820));
sg13g2_nand2_2 U548 (.A(data_o_61_), .B(n904), .Y(n463));
sg13g2_o21ai_1 U550 (.A1(n21), .A2(n905), .B1(n464), .Y(n821));
sg13g2_nand2_2 U551 (.A(data_o_62_), .B(n905), .Y(n464));
sg13g2_o21ai_1 U553 (.A1(n2), .A2(n906), .B1(n465), .Y(n822));
sg13g2_nand2_2 U554 (.A(data_o_63_), .B(n905), .Y(n465));
sg13g2_o21ai_1 U556 (.A1(n356), .A2(n904), .B1(n466), .Y(n823));
sg13g2_nand2_2 U557 (.A(data_o_64_), .B(n904), .Y(n466));
sg13g2_o21ai_1 U559 (.A1(n344), .A2(n907), .B1(n467), .Y(n824));
sg13g2_nand2_2 U560 (.A(data_o_65_), .B(n907), .Y(n467));
sg13g2_o21ai_1 U562 (.A1(n333), .A2(n907), .B1(n468), .Y(n825));
sg13g2_nand2_2 U563 (.A(data_o_66_), .B(n906), .Y(n468));
sg13g2_o21ai_1 U565 (.A1(n322), .A2(n907), .B1(n469), .Y(n826));
sg13g2_nand2_2 U566 (.A(data_o_67_), .B(n904), .Y(n469));
sg13g2_o21ai_1 U568 (.A1(n311), .A2(n906), .B1(n470), .Y(n827));
sg13g2_nand2_2 U569 (.A(data_o_68_), .B(n906), .Y(n470));
sg13g2_o21ai_1 U571 (.A1(n300), .A2(n904), .B1(n471), .Y(n828));
sg13g2_nand2_2 U572 (.A(data_o_69_), .B(n904), .Y(n471));
sg13g2_o21ai_1 U574 (.A1(n289), .A2(n905), .B1(n472), .Y(n829));
sg13g2_nand2_2 U575 (.A(data_o_70_), .B(n904), .Y(n472));
sg13g2_o21ai_1 U577 (.A1(n278), .A2(n906), .B1(n473), .Y(n830));
sg13g2_nand2_2 U578 (.A(data_o_71_), .B(n904), .Y(n473));
sg13g2_o21ai_1 U580 (.A1(n267), .A2(n906), .B1(n474), .Y(n831));
sg13g2_nand2_2 U581 (.A(data_o_72_), .B(n907), .Y(n474));
sg13g2_o21ai_1 U583 (.A1(n256), .A2(n904), .B1(n475), .Y(n832));
sg13g2_nand2_2 U584 (.A(data_o_73_), .B(n907), .Y(n475));
sg13g2_o21ai_1 U586 (.A1(n245), .A2(n904), .B1(n476), .Y(n833));
sg13g2_nand2_2 U587 (.A(data_o_74_), .B(n907), .Y(n476));
sg13g2_o21ai_1 U589 (.A1(n234), .A2(n905), .B1(n477), .Y(n834));
sg13g2_nand2_2 U590 (.A(data_o_75_), .B(n907), .Y(n477));
sg13g2_o21ai_1 U592 (.A1(n223), .A2(n906), .B1(n478), .Y(n835));
sg13g2_nand2_2 U593 (.A(data_o_76_), .B(n904), .Y(n478));
sg13g2_o21ai_1 U595 (.A1(n212), .A2(n906), .B1(n479), .Y(n836));
sg13g2_nand2_2 U596 (.A(data_o_77_), .B(n906), .Y(n479));
sg13g2_o21ai_1 U598 (.A1(n201), .A2(n907), .B1(n480), .Y(n837));
sg13g2_nand2_2 U599 (.A(data_o_78_), .B(n904), .Y(n480));
sg13g2_o21ai_1 U601 (.A1(n190), .A2(n904), .B1(n481), .Y(n838));
sg13g2_nand2_2 U602 (.A(data_o_79_), .B(n907), .Y(n481));
sg13g2_o21ai_1 U604 (.A1(n179), .A2(n906), .B1(n482), .Y(n839));
sg13g2_nand2_2 U605 (.A(data_o_80_), .B(n906), .Y(n482));
sg13g2_o21ai_1 U607 (.A1(n168), .A2(n904), .B1(n483), .Y(n840));
sg13g2_nand2_2 U608 (.A(data_o_81_), .B(n906), .Y(n483));
sg13g2_o21ai_1 U610 (.A1(n157), .A2(n904), .B1(n484), .Y(n841));
sg13g2_nand2_2 U611 (.A(data_o_82_), .B(n904), .Y(n484));
sg13g2_o21ai_1 U613 (.A1(n146), .A2(n906), .B1(n485), .Y(n842));
sg13g2_nand2_2 U614 (.A(data_o_83_), .B(n906), .Y(n485));
sg13g2_o21ai_1 U616 (.A1(n135), .A2(n907), .B1(n486), .Y(n843));
sg13g2_nand2_2 U617 (.A(data_o_84_), .B(n907), .Y(n486));
sg13g2_o21ai_1 U619 (.A1(n124), .A2(n906), .B1(n487), .Y(n844));
sg13g2_nand2_2 U620 (.A(data_o_85_), .B(n904), .Y(n487));
sg13g2_o21ai_1 U622 (.A1(n113), .A2(n904), .B1(n488), .Y(n845));
sg13g2_nand2_2 U623 (.A(data_o_86_), .B(n904), .Y(n488));
sg13g2_o21ai_1 U625 (.A1(n102), .A2(n904), .B1(n489), .Y(n846));
sg13g2_nand2_2 U626 (.A(data_o_87_), .B(n906), .Y(n489));
sg13g2_o21ai_1 U628 (.A1(n91), .A2(n904), .B1(n490), .Y(n847));
sg13g2_nand2_2 U629 (.A(data_o_88_), .B(n906), .Y(n490));
sg13g2_o21ai_1 U631 (.A1(n80), .A2(n905), .B1(n491), .Y(n848));
sg13g2_nand2_2 U632 (.A(data_o_89_), .B(n904), .Y(n491));
sg13g2_o21ai_1 U634 (.A1(n69), .A2(n907), .B1(n492), .Y(n849));
sg13g2_nand2_2 U635 (.A(data_o_90_), .B(n904), .Y(n492));
sg13g2_o21ai_1 U637 (.A1(n58), .A2(n905), .B1(n493), .Y(n850));
sg13g2_nand2_2 U638 (.A(data_o_91_), .B(n904), .Y(n493));
sg13g2_o21ai_1 U640 (.A1(n47), .A2(n907), .B1(n494), .Y(n851));
sg13g2_nand2_2 U641 (.A(data_o_92_), .B(n904), .Y(n494));
sg13g2_o21ai_1 U643 (.A1(n36), .A2(n904), .B1(n495), .Y(n852));
sg13g2_nand2_2 U644 (.A(data_o_93_), .B(n904), .Y(n495));
sg13g2_o21ai_1 U646 (.A1(n25), .A2(n906), .B1(n496), .Y(n853));
sg13g2_nand2_2 U647 (.A(data_o_94_), .B(n905), .Y(n496));
sg13g2_o21ai_1 U649 (.A1(n9), .A2(n907), .B1(n497), .Y(n854));
sg13g2_nand2_2 U650 (.A(data_o_95_), .B(n905), .Y(n497));
sg13g2_o21ai_1 U652 (.A1(n362), .A2(n904), .B1(n498), .Y(n855));
sg13g2_nand2_2 U653 (.A(data_o_96_), .B(n907), .Y(n498));
sg13g2_o21ai_1 U655 (.A1(n348), .A2(n905), .B1(n499), .Y(n856));
sg13g2_nand2_2 U656 (.A(data_o_97_), .B(n905), .Y(n499));
sg13g2_o21ai_1 U658 (.A1(n337), .A2(n904), .B1(n500), .Y(n857));
sg13g2_nand2_2 U659 (.A(data_o_98_), .B(n905), .Y(n500));
sg13g2_o21ai_1 U661 (.A1(n16), .A2(n904), .B1(n501), .Y(n858));
sg13g2_nand2_2 U662 (.A(data_o_127_), .B(n905), .Y(n501));
sg13g2_o21ai_1 U664 (.A1(n29), .A2(n905), .B1(n502), .Y(n859));
sg13g2_nand2_2 U665 (.A(data_o_126_), .B(n907), .Y(n502));
sg13g2_o21ai_1 U667 (.A1(n40), .A2(n907), .B1(n503), .Y(n860));
sg13g2_nand2_2 U668 (.A(data_o_125_), .B(n905), .Y(n503));
sg13g2_o21ai_1 U670 (.A1(n51), .A2(n907), .B1(n504), .Y(n861));
sg13g2_nand2_2 U671 (.A(data_o_124_), .B(n905), .Y(n504));
sg13g2_o21ai_1 U673 (.A1(n62), .A2(n906), .B1(n505), .Y(n862));
sg13g2_nand2_2 U674 (.A(data_o_123_), .B(n906), .Y(n505));
sg13g2_o21ai_1 U676 (.A1(n73), .A2(n906), .B1(n506), .Y(n863));
sg13g2_nand2_2 U677 (.A(data_o_122_), .B(n905), .Y(n506));
sg13g2_o21ai_1 U679 (.A1(n84), .A2(n907), .B1(n507), .Y(n864));
sg13g2_nand2_2 U680 (.A(data_o_121_), .B(n904), .Y(n507));
sg13g2_o21ai_1 U682 (.A1(n95), .A2(n904), .B1(n508), .Y(n865));
sg13g2_nand2_2 U683 (.A(data_o_120_), .B(n904), .Y(n508));
sg13g2_o21ai_1 U685 (.A1(n106), .A2(n907), .B1(n509), .Y(n866));
sg13g2_nand2_2 U686 (.A(data_o_119_), .B(n907), .Y(n509));
sg13g2_o21ai_1 U688 (.A1(n117), .A2(n907), .B1(n510), .Y(n867));
sg13g2_nand2_2 U689 (.A(data_o_118_), .B(n906), .Y(n510));
sg13g2_o21ai_1 U691 (.A1(n128), .A2(n907), .B1(n511), .Y(n868));
sg13g2_nand2_2 U692 (.A(data_o_117_), .B(n907), .Y(n511));
sg13g2_o21ai_1 U694 (.A1(n139), .A2(n906), .B1(n512), .Y(n869));
sg13g2_nand2_2 U695 (.A(data_o_116_), .B(n905), .Y(n512));
sg13g2_o21ai_1 U697 (.A1(n150), .A2(n906), .B1(n513), .Y(n870));
sg13g2_nand2_2 U698 (.A(data_o_115_), .B(n904), .Y(n513));
sg13g2_o21ai_1 U700 (.A1(n161), .A2(n906), .B1(n514), .Y(n871));
sg13g2_nand2_2 U701 (.A(data_o_114_), .B(n905), .Y(n514));
sg13g2_o21ai_1 U703 (.A1(n172), .A2(n907), .B1(n515), .Y(n872));
sg13g2_nand2_2 U704 (.A(data_o_113_), .B(n905), .Y(n515));
sg13g2_o21ai_1 U706 (.A1(n183), .A2(n906), .B1(n516), .Y(n873));
sg13g2_nand2_2 U707 (.A(data_o_112_), .B(n904), .Y(n516));
sg13g2_o21ai_1 U709 (.A1(n194), .A2(n907), .B1(n517), .Y(n874));
sg13g2_nand2_2 U710 (.A(data_o_111_), .B(n905), .Y(n517));
sg13g2_o21ai_1 U712 (.A1(n205), .A2(n907), .B1(n518), .Y(n875));
sg13g2_nand2_2 U713 (.A(data_o_110_), .B(n904), .Y(n518));
sg13g2_o21ai_1 U715 (.A1(n216), .A2(n906), .B1(n519), .Y(n876));
sg13g2_nand2_2 U716 (.A(data_o_109_), .B(n904), .Y(n519));
sg13g2_o21ai_1 U718 (.A1(n227), .A2(n906), .B1(n520), .Y(n877));
sg13g2_nand2_2 U719 (.A(data_o_108_), .B(n904), .Y(n520));
sg13g2_o21ai_1 U721 (.A1(n238), .A2(n907), .B1(n521), .Y(n878));
sg13g2_nand2_2 U722 (.A(data_o_107_), .B(n904), .Y(n521));
sg13g2_o21ai_1 U724 (.A1(n249), .A2(n906), .B1(n522), .Y(n879));
sg13g2_nand2_2 U725 (.A(data_o_106_), .B(n904), .Y(n522));
sg13g2_o21ai_1 U727 (.A1(n260), .A2(n904), .B1(n523), .Y(n880));
sg13g2_nand2_2 U728 (.A(data_o_105_), .B(n904), .Y(n523));
sg13g2_o21ai_1 U730 (.A1(n271), .A2(n906), .B1(n524), .Y(n881));
sg13g2_nand2_2 U731 (.A(data_o_104_), .B(n905), .Y(n524));
sg13g2_o21ai_1 U733 (.A1(n282), .A2(n907), .B1(n525), .Y(n882));
sg13g2_nand2_2 U734 (.A(data_o_103_), .B(n907), .Y(n525));
sg13g2_o21ai_1 U736 (.A1(n293), .A2(n906), .B1(n526), .Y(n883));
sg13g2_nand2_2 U737 (.A(data_o_102_), .B(n906), .Y(n526));
sg13g2_o21ai_1 U739 (.A1(n304), .A2(n907), .B1(n527), .Y(n884));
sg13g2_nand2_2 U740 (.A(data_o_101_), .B(n907), .Y(n527));
sg13g2_o21ai_1 U742 (.A1(n315), .A2(n906), .B1(n528), .Y(n885));
sg13g2_nand2_2 U743 (.A(data_o_100_), .B(n907), .Y(n528));
sg13g2_o21ai_1 U745 (.A1(n326), .A2(n904), .B1(n529), .Y(n886));
sg13g2_nand2_2 U746 (.A(data_o_99_), .B(n906), .Y(n529));
sg13g2_inv_4 U747 (.A(n6), .Y(n896));
sg13g2_inv_4 U748 (.A(n897), .Y(n232));
sg13g2_nand2_2 U750 (.A(n361), .B(n355), .Y(n887));
sg13g2_a21oi_2 U751 (.A1(n355), .A2(n531), .B1(n532), .Y(n888));
sg13g2_nor2_2 U752 (.A(start_i), .B(n531), .Y(n532));
sg13g2_nand2_2 U753 (.A(outy_20_), .B(n896), .Y(n898));
sg13g2_nand2_2 U754 (.A(data_i_41_), .B(n1), .Y(n536));
sg13g2_nand2_2 U755 (.A(data_i_73_), .B(n8), .Y(n535));
sg13g2_nand2_2 U756 (.A(data_i_105_), .B(n15), .Y(n534));
sg13g2_nand2_2 U757 (.A(data_i_9_), .B(next_ready_o), .Y(n533));
sg13g2_inv_4 U758 (.A(n898), .Y(n133));
sg13g2_nand2_2 U759 (.A(data_i_40_), .B(n1), .Y(n540));
sg13g2_nand2_2 U760 (.A(data_i_72_), .B(n8), .Y(n539));
sg13g2_nand2_2 U761 (.A(data_i_104_), .B(n15), .Y(n538));
sg13g2_nand2_2 U762 (.A(data_i_8_), .B(next_ready_o), .Y(n537));
sg13g2_o21ai_1 U763 (.A1(n1), .A2(n219), .B1(n220), .Y(n720));
sg13g2_nand2_2 U764 (.A(data_i_53_), .B(n1), .Y(n608));
sg13g2_nand2_2 U765 (.A(data_i_127_), .B(n15), .Y(n562));
sg13g2_nand2_2 U766 (.A(data_i_103_), .B(n15), .Y(n542));
sg13g2_nand2_2 U767 (.A(data_i_7_), .B(next_ready_o), .Y(n541));
sg13g2_o21ai_1 U768 (.A1(n1), .A2(n109), .B1(n110), .Y(n690));
sg13g2_nand2_2 U769 (.A(data_i_38_), .B(n1), .Y(n548));
sg13g2_nand2_2 U770 (.A(data_i_70_), .B(n8), .Y(n547));
sg13g2_nand2_2 U771 (.A(data_i_102_), .B(n15), .Y(n546));
sg13g2_nand2_2 U772 (.A(data_i_6_), .B(next_ready_o), .Y(n545));
sg13g2_nor2_2 U773 (.A(n112), .B(n6), .Y(n111));
sg13g2_nand2_2 U774 (.A(data_i_37_), .B(n1), .Y(n552));
sg13g2_nand2_2 U775 (.A(data_i_69_), .B(n8), .Y(n551));
sg13g2_nand2_2 U776 (.A(data_i_101_), .B(n15), .Y(n550));
sg13g2_nand2_2 U777 (.A(data_i_5_), .B(next_ready_o), .Y(n549));
sg13g2_nand2_2 U778 (.A(data_i_45_), .B(n1), .Y(n644));
sg13g2_nand2_2 U779 (.A(data_i_36_), .B(n1), .Y(n556));
sg13g2_nand2_2 U780 (.A(data_i_68_), .B(n8), .Y(n555));
sg13g2_nand2_2 U781 (.A(data_i_100_), .B(n15), .Y(n554));
sg13g2_nand2_2 U782 (.A(data_i_4_), .B(next_ready_o), .Y(n553));
sg13g2_nand2_2 U783 (.A(data_i_61_), .B(n1), .Y(n576));
sg13g2_nand2_2 U784 (.A(data_i_35_), .B(n1), .Y(n560));
sg13g2_nand2_2 U785 (.A(data_i_67_), .B(n8), .Y(n559));
sg13g2_nand2_2 U786 (.A(data_i_99_), .B(n15), .Y(n558));
sg13g2_nand2_2 U787 (.A(data_i_3_), .B(next_ready_o), .Y(n557));
sg13g2_nand2_2 U788 (.A(data_i_125_), .B(n15), .Y(n574));
sg13g2_nand4_1 U789 (.A(n545), .B(n546), .C(n547), .D(n548), .Y(mix_word_6_));
sg13g2_nand2_2 U790 (.A(data_i_95_), .B(n8), .Y(n563));
sg13g2_nand4_1 U791 (.A(n577), .B(n578), .C(n579), .D(n580), .Y(mix_word_28_));
sg13g2_nand2_2 U792 (.A(data_i_31_), .B(next_ready_o), .Y(n561));
sg13g2_nor2_2 U793 (.A(n20), .B(n226), .Y(n229));
sg13g2_nand4_1 U794 (.A(n609), .B(n610), .C(n611), .D(n612), .Y(mix_word_20_));
sg13g2_nand2_2 U795 (.A(data_i_94_), .B(n8), .Y(n567));
sg13g2_nand2_2 U796 (.A(data_i_126_), .B(n15), .Y(n566));
sg13g2_nand2_2 U797 (.A(data_i_30_), .B(next_ready_o), .Y(n565));
sg13g2_o21ai_1 U798 (.A1(n15), .A2(n139), .B1(n140), .Y(n698));
sg13g2_nand2_2 U799 (.A(data_i_34_), .B(n1), .Y(n572));
sg13g2_nand2_2 U800 (.A(data_i_66_), .B(n8), .Y(n571));
sg13g2_nand2_2 U801 (.A(data_i_98_), .B(n15), .Y(n570));
sg13g2_nand2_2 U802 (.A(data_i_2_), .B(next_ready_o), .Y(n569));
sg13g2_nand4_1 U803 (.A(n645), .B(n646), .C(n647), .D(n648), .Y(mix_word_12_));
sg13g2_o21ai_1 U804 (.A1(n15), .A2(n315), .B1(n316), .Y(n746));
sg13g2_o21ai_1 U805 (.A1(n8), .A2(n135), .B1(n136), .Y(n697));
sg13g2_o21ai_1 U806 (.A1(n8), .A2(n311), .B1(n312), .Y(n745));
sg13g2_nand2_2 U807 (.A(data_i_29_), .B(next_ready_o), .Y(n573));
sg13g2_o21ai_1 U808 (.A1(n8), .A2(n223), .B1(n224), .Y(n721));
sg13g2_nand2_2 U809 (.A(data_i_60_), .B(n1), .Y(n580));
sg13g2_nand2_2 U810 (.A(data_i_92_), .B(n8), .Y(n579));
sg13g2_nand2_2 U811 (.A(data_i_124_), .B(n15), .Y(n578));
sg13g2_nand2_2 U812 (.A(data_i_28_), .B(next_ready_o), .Y(n577));
sg13g2_nand4_1 U813 (.A(n553), .B(n554), .C(n555), .D(n556), .Y(mix_word_4_));
sg13g2_nand2_2 U814 (.A(data_i_59_), .B(n1), .Y(n584));
sg13g2_nand2_2 U815 (.A(data_i_91_), .B(n8), .Y(n583));
sg13g2_nand2_2 U816 (.A(data_i_123_), .B(n15), .Y(n582));
sg13g2_nand2_2 U817 (.A(data_i_27_), .B(next_ready_o), .Y(n581));
sg13g2_nor2_2 U818 (.A(n899), .B(n369), .Y(n900));
sg13g2_nand2_2 U819 (.A(data_i_58_), .B(n1), .Y(n588));
sg13g2_nand2_2 U820 (.A(data_i_90_), .B(n8), .Y(n587));
sg13g2_nand2_2 U821 (.A(data_i_122_), .B(n15), .Y(n586));
sg13g2_nand2_2 U822 (.A(data_i_26_), .B(next_ready_o), .Y(n585));
sg13g2_inv_4 U823 (.A(outx_19_), .Y(n899));
sg13g2_nand2_2 U824 (.A(data_i_57_), .B(n1), .Y(n592));
sg13g2_nand2_2 U825 (.A(data_i_89_), .B(n8), .Y(n591));
sg13g2_nand2_2 U826 (.A(data_i_121_), .B(n15), .Y(n590));
sg13g2_nand2_2 U827 (.A(data_i_25_), .B(next_ready_o), .Y(n589));
sg13g2_o21ai_1 U828 (.A1(n1), .A2(n318), .B1(n319), .Y(n747));
sg13g2_nand2_2 U829 (.A(data_i_56_), .B(n1), .Y(n596));
sg13g2_nand2_2 U830 (.A(data_i_88_), .B(n8), .Y(n595));
sg13g2_nand2_2 U831 (.A(data_i_120_), .B(n15), .Y(n594));
sg13g2_nand2_2 U832 (.A(data_i_24_), .B(next_ready_o), .Y(n593));
sg13g2_o21ai_1 U833 (.A1(n1), .A2(n120), .B1(n121), .Y(n693));
sg13g2_nand2_2 U834 (.A(data_i_55_), .B(n1), .Y(n600));
sg13g2_nand2_2 U835 (.A(data_i_87_), .B(n8), .Y(n599));
sg13g2_nand2_2 U836 (.A(data_i_119_), .B(n15), .Y(n598));
sg13g2_nand2_2 U837 (.A(data_i_23_), .B(next_ready_o), .Y(n597));
sg13g2_nand2_2 U838 (.A(n355), .B(data_reg_62_), .Y(n901));
sg13g2_nand2_2 U839 (.A(data_i_54_), .B(n1), .Y(n604));
sg13g2_nand2_2 U840 (.A(data_i_86_), .B(n8), .Y(n603));
sg13g2_nand2_2 U841 (.A(data_i_118_), .B(n15), .Y(n602));
sg13g2_nand2_2 U842 (.A(data_i_22_), .B(next_ready_o), .Y(n601));
sg13g2_inv_4 U843 (.A(outx_30_), .Y(n902));
sg13g2_nor2_2 U844 (.A(n6), .B(n892), .Y(n298));
sg13g2_nand2_2 U845 (.A(data_i_62_), .B(n1), .Y(n568));
sg13g2_nand4_1 U846 (.A(n629), .B(n630), .C(n631), .D(n632), .Y(mix_word_16_));
sg13g2_nand2_2 U847 (.A(data_i_77_), .B(n8), .Y(n643));
sg13g2_nand4_1 U848 (.A(n625), .B(n626), .C(n627), .D(n628), .Y(mix_word_17_));
sg13g2_nand2_2 U849 (.A(data_i_52_), .B(n1), .Y(n612));
sg13g2_nand2_2 U850 (.A(data_i_84_), .B(n8), .Y(n611));
sg13g2_nand2_2 U851 (.A(data_i_116_), .B(n15), .Y(n610));
sg13g2_nand2_2 U852 (.A(data_i_20_), .B(next_ready_o), .Y(n609));
sg13g2_nand4_1 U853 (.A(n589), .B(n590), .C(n591), .D(n592), .Y(mix_word_25_));
sg13g2_nand2_2 U854 (.A(data_i_33_), .B(n1), .Y(n616));
sg13g2_nand2_2 U855 (.A(data_i_65_), .B(n8), .Y(n615));
sg13g2_nand2_2 U856 (.A(data_i_97_), .B(n15), .Y(n614));
sg13g2_nand2_2 U857 (.A(data_i_1_), .B(next_ready_o), .Y(n613));
sg13g2_o21ai_1 U858 (.A1(n1), .A2(n175), .B1(n176), .Y(n708));
sg13g2_nand2_2 U859 (.A(data_i_51_), .B(n1), .Y(n620));
sg13g2_nand2_2 U860 (.A(data_i_83_), .B(n8), .Y(n619));
sg13g2_nand2_2 U861 (.A(data_i_115_), .B(n15), .Y(n618));
sg13g2_nand2_2 U862 (.A(data_i_19_), .B(next_ready_o), .Y(n617));
sg13g2_o21ai_1 U863 (.A1(n1), .A2(n263), .B1(n264), .Y(n732));
sg13g2_nand2_2 U864 (.A(data_i_50_), .B(n1), .Y(n624));
sg13g2_nand2_2 U865 (.A(data_i_82_), .B(n8), .Y(n623));
sg13g2_nand2_2 U866 (.A(data_i_114_), .B(n15), .Y(n622));
sg13g2_nand2_2 U867 (.A(data_i_18_), .B(next_ready_o), .Y(n621));
sg13g2_nand4_1 U868 (.A(n533), .B(n534), .C(n535), .D(n536), .Y(mix_word_9_));
sg13g2_nand2_2 U869 (.A(data_i_49_), .B(n1), .Y(n628));
sg13g2_nand2_2 U870 (.A(data_i_81_), .B(n8), .Y(n627));
sg13g2_nand2_2 U871 (.A(data_i_113_), .B(n15), .Y(n626));
sg13g2_nand2_2 U872 (.A(data_i_17_), .B(next_ready_o), .Y(n625));
sg13g2_nor2_2 U873 (.A(n6), .B(n321), .Y(n320));
sg13g2_nand2_2 U874 (.A(data_i_48_), .B(n1), .Y(n632));
sg13g2_nand2_2 U875 (.A(data_i_80_), .B(n8), .Y(n631));
sg13g2_nand2_2 U876 (.A(data_i_112_), .B(n15), .Y(n630));
sg13g2_nand2_2 U877 (.A(data_i_16_), .B(next_ready_o), .Y(n629));
sg13g2_o21ai_1 U878 (.A1(n1), .A2(n208), .B1(n209), .Y(n717));
sg13g2_nand2_2 U879 (.A(data_i_47_), .B(n1), .Y(n636));
sg13g2_nand2_2 U880 (.A(data_i_79_), .B(n8), .Y(n635));
sg13g2_nand2_2 U881 (.A(data_i_111_), .B(n15), .Y(n634));
sg13g2_nand2_2 U882 (.A(data_i_15_), .B(next_ready_o), .Y(n633));
sg13g2_o21ai_1 U883 (.A1(n15), .A2(n84), .B1(n85), .Y(n683));
sg13g2_nand2_2 U884 (.A(data_i_46_), .B(n1), .Y(n640));
sg13g2_nand2_2 U885 (.A(data_i_78_), .B(n8), .Y(n639));
sg13g2_nand2_2 U886 (.A(data_i_110_), .B(n15), .Y(n638));
sg13g2_nand2_2 U887 (.A(data_i_14_), .B(next_ready_o), .Y(n637));
sg13g2_o21ai_1 U888 (.A1(n8), .A2(n80), .B1(n81), .Y(n682));
sg13g2_nand4_1 U889 (.A(n653), .B(n654), .C(n655), .D(n656), .Y(mix_word_10_));
sg13g2_nand4_1 U890 (.A(n585), .B(n586), .C(n587), .D(n588), .Y(mix_word_26_));
sg13g2_nand4_1 U891 (.A(n569), .B(n570), .C(n571), .D(n572), .Y(mix_word_2_));
sg13g2_nor2_2 U892 (.A(n6), .B(n890), .Y(n309));
sg13g2_nand4_1 U893 (.A(n621), .B(n622), .C(n623), .D(n624), .Y(mix_word_18_));
sg13g2_nand2_2 U894 (.A(data_i_44_), .B(n1), .Y(n648));
sg13g2_nand2_2 U895 (.A(data_i_76_), .B(n8), .Y(n647));
sg13g2_nand2_2 U896 (.A(data_i_108_), .B(n15), .Y(n646));
sg13g2_nand2_2 U897 (.A(data_i_12_), .B(next_ready_o), .Y(n645));
sg13g2_nand4_1 U898 (.A(n613), .B(n614), .C(n615), .D(n616), .Y(mix_word_1_));
sg13g2_nand2_2 U899 (.A(data_i_43_), .B(n1), .Y(n652));
sg13g2_nand2_2 U900 (.A(data_i_75_), .B(n8), .Y(n651));
sg13g2_nand2_2 U901 (.A(data_i_107_), .B(n15), .Y(n650));
sg13g2_nand2_2 U902 (.A(data_i_11_), .B(next_ready_o), .Y(n649));
sg13g2_nand4_1 U903 (.A(n617), .B(n618), .C(n619), .D(n620), .Y(mix_word_19_));
sg13g2_nand2_2 U904 (.A(data_i_42_), .B(n1), .Y(n656));
sg13g2_nand2_2 U905 (.A(data_i_74_), .B(n8), .Y(n655));
sg13g2_nand2_2 U906 (.A(data_i_106_), .B(n15), .Y(n654));
sg13g2_nand2_2 U907 (.A(data_i_10_), .B(next_ready_o), .Y(n653));
sg13g2_nand4_1 U908 (.A(n581), .B(n582), .C(n583), .D(n584), .Y(mix_word_27_));
sg13g2_nand2_2 U909 (.A(data_i_32_), .B(n1), .Y(n660));
sg13g2_nand4_1 U910 (.A(n649), .B(n650), .C(n651), .D(n652), .Y(mix_word_11_));
sg13g2_nor2_2 U911 (.A(n6), .B(n24), .Y(n23));
sg13g2_nand2_2 U912 (.A(data_i_64_), .B(n8), .Y(n659));
sg13g2_nand4_1 U913 (.A(n557), .B(n558), .C(n559), .D(n560), .Y(mix_word_3_));
sg13g2_nor2_2 U914 (.A(n6), .B(n288), .Y(n287));
sg13g2_nand2_2 U915 (.A(data_i_96_), .B(n15), .Y(n658));
sg13g2_o21ai_1 U916 (.A1(n1), .A2(n351), .B1(n352), .Y(n756));
sg13g2_nor2_2 U917 (.A(n6), .B(n90), .Y(n89));
sg13g2_inv_4 U918 (.A(n531), .Y(n530));
sg13g2_nand2_2 U919 (.A(n661), .B(n662), .Y(n531));
sg13g2_nand2_2 U920 (.A(data_i_0_), .B(next_ready_o), .Y(n657));
sg13g2_nand4_1 U921 (.A(n537), .B(n538), .C(n539), .D(n540), .Y(mix_word_8_));
sg13g2_nand4_1 U922 (.A(n657), .B(n658), .C(n659), .D(n660), .Y(mix_word_0_));
sg13g2_nand4_1 U923 (.A(n633), .B(n634), .C(n635), .D(n636), .Y(mix_word_15_));
sg13g2_nand4_1 U924 (.A(n541), .B(n542), .C(n543), .D(n544), .Y(mix_word_7_));
sg13g2_nand4_1 U925 (.A(n597), .B(n598), .C(n599), .D(n600), .Y(mix_word_23_));
sg13g2_o21ai_1 U926 (.A1(n1), .A2(n54), .B1(n55), .Y(n675));
sg13g2_o21ai_1 U927 (.A1(n1), .A2(n131), .B1(n132), .Y(n696));
sg13g2_nand4_1 U928 (.A(n561), .B(n562), .C(n563), .D(n564), .Y(mix_word_31_));
sg13g2_nand4_1 U929 (.A(n641), .B(n642), .C(n643), .D(n644), .Y(mix_word_13_));
sg13g2_nand4_1 U930 (.A(n565), .B(n566), .C(n567), .D(n568), .Y(mix_word_30_));
sg13g2_inv_4 U931 (.A(n361), .Y(n8));
sg13g2_nand4_1 U932 (.A(n607), .B(n606), .C(n605), .D(n608), .Y(mix_word_21_));
sg13g2_inv_4 U933 (.A(n355), .Y(n1));
sg13g2_nand4_1 U934 (.A(n552), .B(n550), .C(n551), .D(n549), .Y(mix_word_5_));
sg13g2_o21ai_1 U935 (.A1(n1), .A2(n43), .B1(n44), .Y(n672));
sg13g2_nand4_1 U936 (.A(n601), .B(n602), .C(n603), .D(n604), .Y(mix_word_22_));
sg13g2_inv_4 U937 (.A(n365), .Y(n15));
sg13g2_nand2_2 U938 (.A(start_i), .B(n530), .Y(n365));
sg13g2_inv_4 U939 (.A(n433), .Y(n904));
sg13g2_inv_4 U940 (.A(n433), .Y(n907));
sg13g2_inv_4 U941 (.A(n433), .Y(n905));
sg13g2_inv_4 U942 (.A(n433), .Y(n906));
sg13g2_dfrbp_1 data_o_reg_reg_0_ (.CLK(clk), .D(n759), .Q(data_o_0_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_1_ (.CLK(clk), .D(n760), .Q(data_o_1_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_2_ (.CLK(clk), .D(n761), .Q(data_o_2_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_3_ (.CLK(clk), .D(n762), .Q(data_o_3_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_4_ (.CLK(clk), .D(n763), .Q(data_o_4_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_5_ (.CLK(clk), .D(n764), .Q(data_o_5_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_6_ (.CLK(clk), .D(n765), .Q(data_o_6_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_7_ (.CLK(clk), .D(n766), .Q(data_o_7_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_8_ (.CLK(clk), .D(n767), .Q(data_o_8_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_9_ (.CLK(clk), .D(n768), .Q(data_o_9_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_10_ (.CLK(clk), .D(n769), .Q(data_o_10_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_11_ (.CLK(clk), .D(n770), .Q(data_o_11_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_12_ (.CLK(clk), .D(n771), .Q(data_o_12_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_13_ (.CLK(clk), .D(n772), .Q(data_o_13_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_14_ (.CLK(clk), .D(n773), .Q(data_o_14_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_15_ (.CLK(clk), .D(n774), .Q(data_o_15_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_16_ (.CLK(clk), .D(n775), .Q(data_o_16_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_17_ (.CLK(clk), .D(n776), .Q(data_o_17_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_18_ (.CLK(clk), .D(n777), .Q(data_o_18_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_19_ (.CLK(clk), .D(n778), .Q(data_o_19_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_20_ (.CLK(clk), .D(n779), .Q(data_o_20_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_21_ (.CLK(clk), .D(n780), .Q(data_o_21_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_22_ (.CLK(clk), .D(n781), .Q(data_o_22_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_23_ (.CLK(clk), .D(n782), .Q(data_o_23_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_24_ (.CLK(clk), .D(n783), .Q(data_o_24_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_25_ (.CLK(clk), .D(n784), .Q(data_o_25_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_26_ (.CLK(clk), .D(n785), .Q(data_o_26_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_27_ (.CLK(clk), .D(n786), .Q(data_o_27_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_28_ (.CLK(clk), .D(n787), .Q(data_o_28_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_29_ (.CLK(clk), .D(n788), .Q(data_o_29_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_30_ (.CLK(clk), .D(n789), .Q(data_o_30_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_31_ (.CLK(clk), .D(n790), .Q(data_o_31_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_32_ (.CLK(clk), .D(n791), .Q(data_o_32_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_33_ (.CLK(clk), .D(n792), .Q(data_o_33_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_34_ (.CLK(clk), .D(n793), .Q(data_o_34_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_35_ (.CLK(clk), .D(n794), .Q(data_o_35_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_36_ (.CLK(clk), .D(n795), .Q(data_o_36_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_37_ (.CLK(clk), .D(n796), .Q(data_o_37_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_38_ (.CLK(clk), .D(n797), .Q(data_o_38_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_39_ (.CLK(clk), .D(n798), .Q(data_o_39_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_40_ (.CLK(clk), .D(n799), .Q(data_o_40_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_41_ (.CLK(clk), .D(n800), .Q(data_o_41_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_42_ (.CLK(clk), .D(n801), .Q(data_o_42_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_43_ (.CLK(clk), .D(n802), .Q(data_o_43_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_44_ (.CLK(clk), .D(n803), .Q(data_o_44_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_45_ (.CLK(clk), .D(n804), .Q(data_o_45_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_46_ (.CLK(clk), .D(n805), .Q(data_o_46_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_47_ (.CLK(clk), .D(n806), .Q(data_o_47_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_48_ (.CLK(clk), .D(n807), .Q(data_o_48_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_49_ (.CLK(clk), .D(n808), .Q(data_o_49_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_50_ (.CLK(clk), .D(n809), .Q(data_o_50_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_51_ (.CLK(clk), .D(n810), .Q(data_o_51_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_52_ (.CLK(clk), .D(n811), .Q(data_o_52_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_53_ (.CLK(clk), .D(n812), .Q(data_o_53_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_54_ (.CLK(clk), .D(n813), .Q(data_o_54_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_55_ (.CLK(clk), .D(n814), .Q(data_o_55_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_56_ (.CLK(clk), .D(n815), .Q(data_o_56_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_57_ (.CLK(clk), .D(n816), .Q(data_o_57_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_58_ (.CLK(clk), .D(n817), .Q(data_o_58_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_59_ (.CLK(clk), .D(n818), .Q(data_o_59_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_60_ (.CLK(clk), .D(n819), .Q(data_o_60_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_61_ (.CLK(clk), .D(n820), .Q(data_o_61_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_62_ (.CLK(clk), .D(n821), .Q(data_o_62_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_63_ (.CLK(clk), .D(n822), .Q(data_o_63_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_64_ (.CLK(clk), .D(n823), .Q(data_o_64_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_65_ (.CLK(clk), .D(n824), .Q(data_o_65_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_66_ (.CLK(clk), .D(n825), .Q(data_o_66_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_67_ (.CLK(clk), .D(n826), .Q(data_o_67_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_68_ (.CLK(clk), .D(n827), .Q(data_o_68_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_69_ (.CLK(clk), .D(n828), .Q(data_o_69_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_70_ (.CLK(clk), .D(n829), .Q(data_o_70_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_71_ (.CLK(clk), .D(n830), .Q(data_o_71_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_72_ (.CLK(clk), .D(n831), .Q(data_o_72_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_73_ (.CLK(clk), .D(n832), .Q(data_o_73_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_74_ (.CLK(clk), .D(n833), .Q(data_o_74_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_75_ (.CLK(clk), .D(n834), .Q(data_o_75_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_76_ (.CLK(clk), .D(n835), .Q(data_o_76_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_77_ (.CLK(clk), .D(n836), .Q(data_o_77_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_78_ (.CLK(clk), .D(n837), .Q(data_o_78_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_79_ (.CLK(clk), .D(n838), .Q(data_o_79_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_80_ (.CLK(clk), .D(n839), .Q(data_o_80_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_81_ (.CLK(clk), .D(n840), .Q(data_o_81_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_82_ (.CLK(clk), .D(n841), .Q(data_o_82_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_83_ (.CLK(clk), .D(n842), .Q(data_o_83_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_84_ (.CLK(clk), .D(n843), .Q(data_o_84_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_85_ (.CLK(clk), .D(n844), .Q(data_o_85_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_86_ (.CLK(clk), .D(n845), .Q(data_o_86_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_87_ (.CLK(clk), .D(n846), .Q(data_o_87_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_88_ (.CLK(clk), .D(n847), .Q(data_o_88_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_89_ (.CLK(clk), .D(n848), .Q(data_o_89_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_90_ (.CLK(clk), .D(n849), .Q(data_o_90_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_91_ (.CLK(clk), .D(n850), .Q(data_o_91_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_92_ (.CLK(clk), .D(n851), .Q(data_o_92_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_93_ (.CLK(clk), .D(n852), .Q(data_o_93_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_94_ (.CLK(clk), .D(n853), .Q(data_o_94_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_95_ (.CLK(clk), .D(n854), .Q(data_o_95_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_96_ (.CLK(clk), .D(n855), .Q(data_o_96_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_97_ (.CLK(clk), .D(n856), .Q(data_o_97_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_98_ (.CLK(clk), .D(n857), .Q(data_o_98_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_99_ (.CLK(clk), .D(n886), .Q(data_o_99_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_100_ (.CLK(clk), .D(n885), .Q(data_o_100_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_101_ (.CLK(clk), .D(n884), .Q(data_o_101_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_102_ (.CLK(clk), .D(n883), .Q(data_o_102_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_103_ (.CLK(clk), .D(n882), .Q(data_o_103_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_104_ (.CLK(clk), .D(n881), .Q(data_o_104_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_105_ (.CLK(clk), .D(n880), .Q(data_o_105_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_106_ (.CLK(clk), .D(n879), .Q(data_o_106_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_107_ (.CLK(clk), .D(n878), .Q(data_o_107_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_108_ (.CLK(clk), .D(n877), .Q(data_o_108_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_109_ (.CLK(clk), .D(n876), .Q(data_o_109_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_110_ (.CLK(clk), .D(n875), .Q(data_o_110_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_111_ (.CLK(clk), .D(n874), .Q(data_o_111_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_112_ (.CLK(clk), .D(n873), .Q(data_o_112_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_113_ (.CLK(clk), .D(n872), .Q(data_o_113_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_114_ (.CLK(clk), .D(n871), .Q(data_o_114_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_115_ (.CLK(clk), .D(n870), .Q(data_o_115_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_116_ (.CLK(clk), .D(n869), .Q(data_o_116_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_117_ (.CLK(clk), .D(n868), .Q(data_o_117_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_118_ (.CLK(clk), .D(n867), .Q(data_o_118_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_119_ (.CLK(clk), .D(n866), .Q(data_o_119_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_120_ (.CLK(clk), .D(n865), .Q(data_o_120_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_121_ (.CLK(clk), .D(n864), .Q(data_o_121_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_122_ (.CLK(clk), .D(n863), .Q(data_o_122_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_123_ (.CLK(clk), .D(n862), .Q(data_o_123_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_124_ (.CLK(clk), .D(n861), .Q(data_o_124_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_125_ (.CLK(clk), .D(n860), .Q(data_o_125_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_126_ (.CLK(clk), .D(n859), .Q(data_o_126_), .RESET_B(reset));
sg13g2_dfrbp_1 data_o_reg_reg_127_ (.CLK(clk), .D(n858), .Q(data_o_127_), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_32_ (.CLK(clk), .D(n756), .Q_N(n351), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_33_ (.CLK(clk), .D(n753), .Q_N(n340), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_34_ (.CLK(clk), .D(n750), .Q_N(n329), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_35_ (.CLK(clk), .D(n747), .Q_N(n318), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_36_ (.CLK(clk), .D(n744), .Q_N(n307), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_37_ (.CLK(clk), .D(n741), .Q_N(n296), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_38_ (.CLK(clk), .D(n738), .Q_N(n285), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_39_ (.CLK(clk), .D(n735), .Q_N(n274), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_40_ (.CLK(clk), .D(n732), .Q_N(n263), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_41_ (.CLK(clk), .D(n729), .Q_N(n252), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_42_ (.CLK(clk), .D(n726), .Q_N(n241), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_43_ (.CLK(clk), .D(n723), .Q_N(n230), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_44_ (.CLK(clk), .D(n720), .Q_N(n219), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_45_ (.CLK(clk), .D(n717), .Q_N(n208), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_46_ (.CLK(clk), .D(n714), .Q_N(n197), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_47_ (.CLK(clk), .D(n711), .Q_N(n186), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_48_ (.CLK(clk), .D(n708), .Q_N(n175), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_49_ (.CLK(clk), .D(n705), .Q_N(n164), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_50_ (.CLK(clk), .D(n702), .Q_N(n153), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_51_ (.CLK(clk), .D(n699), .Q_N(n142), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_52_ (.CLK(clk), .D(n696), .Q_N(n131), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_53_ (.CLK(clk), .D(n693), .Q_N(n120), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_54_ (.CLK(clk), .D(n690), .Q_N(n109), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_55_ (.CLK(clk), .D(n687), .Q_N(n98), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_56_ (.CLK(clk), .D(n684), .Q_N(n87), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_57_ (.CLK(clk), .D(n681), .Q_N(n76), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_58_ (.CLK(clk), .D(n678), .Q_N(n65), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_59_ (.CLK(clk), .D(n675), .Q_N(n54), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_60_ (.CLK(clk), .D(n672), .Q_N(n43), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_61_ (.CLK(clk), .D(n669), .Q_N(n32), .RESET_B(reset));
sg13g2_dfrbp_1 data_reg_reg_62_ (.CLK(clk), .D(n666), .Q(data_reg_62_), .Q_N(n21), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_63_ (.CLK(clk), .D(n663), .Q_N(n2), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_64_ (.CLK(clk), .D(n757), .Q_N(n356), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_65_ (.CLK(clk), .D(n754), .Q_N(n344), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_66_ (.CLK(clk), .D(n751), .Q_N(n333), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_67_ (.CLK(clk), .D(n748), .Q_N(n322), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_68_ (.CLK(clk), .D(n745), .Q_N(n311), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_69_ (.CLK(clk), .D(n742), .Q_N(n300), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_70_ (.CLK(clk), .D(n739), .Q_N(n289), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_71_ (.CLK(clk), .D(n736), .Q_N(n278), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_72_ (.CLK(clk), .D(n733), .Q_N(n267), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_73_ (.CLK(clk), .D(n730), .Q_N(n256), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_74_ (.CLK(clk), .D(n727), .Q_N(n245), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_75_ (.CLK(clk), .D(n724), .Q_N(n234), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_76_ (.CLK(clk), .D(n721), .Q_N(n223), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_77_ (.CLK(clk), .D(n718), .Q_N(n212), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_78_ (.CLK(clk), .D(n715), .Q_N(n201), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_79_ (.CLK(clk), .D(n712), .Q_N(n190), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_80_ (.CLK(clk), .D(n709), .Q_N(n179), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_81_ (.CLK(clk), .D(n706), .Q_N(n168), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_82_ (.CLK(clk), .D(n703), .Q_N(n157), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_83_ (.CLK(clk), .D(n700), .Q_N(n146), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_84_ (.CLK(clk), .D(n697), .Q_N(n135), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_85_ (.CLK(clk), .D(n694), .Q_N(n124), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_86_ (.CLK(clk), .D(n691), .Q_N(n113), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_87_ (.CLK(clk), .D(n688), .Q_N(n102), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_88_ (.CLK(clk), .D(n685), .Q_N(n91), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_89_ (.CLK(clk), .D(n682), .Q_N(n80), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_90_ (.CLK(clk), .D(n679), .Q_N(n69), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_91_ (.CLK(clk), .D(n676), .Q_N(n58), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_92_ (.CLK(clk), .D(n673), .Q_N(n47), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_93_ (.CLK(clk), .D(n670), .Q_N(n36), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_94_ (.CLK(clk), .D(n667), .Q_N(n25), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_95_ (.CLK(clk), .D(n664), .Q_N(n9), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_96_ (.CLK(clk), .D(n758), .Q_N(n362), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_97_ (.CLK(clk), .D(n755), .Q_N(n348), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_98_ (.CLK(clk), .D(n752), .Q_N(n337), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_99_ (.CLK(clk), .D(n749), .Q_N(n326), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_100_ (.CLK(clk), .D(n746), .Q_N(n315), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_101_ (.CLK(clk), .D(n743), .Q_N(n304), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_102_ (.CLK(clk), .D(n740), .Q_N(n293), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_103_ (.CLK(clk), .D(n737), .Q_N(n282), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_104_ (.CLK(clk), .D(n734), .Q_N(n271), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_105_ (.CLK(clk), .D(n731), .Q_N(n260), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_106_ (.CLK(clk), .D(n728), .Q_N(n249), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_107_ (.CLK(clk), .D(n725), .Q_N(n238), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_108_ (.CLK(clk), .D(n722), .Q_N(n227), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_109_ (.CLK(clk), .D(n719), .Q_N(n216), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_110_ (.CLK(clk), .D(n716), .Q_N(n205), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_111_ (.CLK(clk), .D(n713), .Q_N(n194), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_112_ (.CLK(clk), .D(n710), .Q_N(n183), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_113_ (.CLK(clk), .D(n707), .Q_N(n172), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_114_ (.CLK(clk), .D(n704), .Q_N(n161), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_115_ (.CLK(clk), .D(n701), .Q_N(n150), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_116_ (.CLK(clk), .D(n698), .Q_N(n139), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_117_ (.CLK(clk), .D(n695), .Q_N(n128), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_118_ (.CLK(clk), .D(n692), .Q_N(n117), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_119_ (.CLK(clk), .D(n689), .Q_N(n106), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_120_ (.CLK(clk), .D(n686), .Q_N(n95), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_121_ (.CLK(clk), .D(n683), .Q_N(n84), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_122_ (.CLK(clk), .D(n680), .Q_N(n73), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_123_ (.CLK(clk), .D(n677), .Q_N(n62), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_124_ (.CLK(clk), .D(n674), .Q_N(n51), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_125_ (.CLK(clk), .D(n671), .Q_N(n40), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_126_ (.CLK(clk), .D(n668), .Q_N(n29), .RESET_B(reset));
sg13g2_dfrbp_2 data_reg_reg_127_ (.CLK(clk), .D(n665), .Q_N(n16), .RESET_B(reset));
sg13g2_dfrbp_1 ready_o_reg (.CLK(clk), .D(next_ready_o), .Q(ready_o), .RESET_B(reset));
sg13g2_dfrbp_2 state_reg_0_ (.CLK(clk), .D(n888), .Q(state_0_), .Q_N(n661), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_1_ (.CLK(clk), .D(n887), .Q(state_1_), .Q_N(n662), .RESET_B(reset));
word_mixcolum w1(.in_0_(mix_word_0_), .in_1_(mix_word_1_), .in_2_(mix_word_2_), .in_3_(mix_word_3_), .in_4_(mix_word_4_), .in_5_(mix_word_5_), .in_6_(mix_word_6_), .in_7_(mix_word_7_), .in_8_(mix_word_8_), .in_9_(mix_word_9_), .in_10_(mix_word_10_), .in_11_(mix_word_11_), .in_12_(mix_word_12_), .in_13_(mix_word_13_), .in_14_(mix_word_14_), .in_15_(mix_word_15_), .in_16_(mix_word_16_), .in_17_(mix_word_17_), .in_18_(mix_word_18_), .in_19_(mix_word_19_), .in_20_(mix_word_20_), .in_21_(mix_word_21_), .in_22_(mix_word_22_), .in_23_(mix_word_23_), .in_24_(mix_word_24_), .in_25_(mix_word_25_), .in_26_(mix_word_26_), .in_27_(mix_word_27_), .in_28_(mix_word_28_), .in_29_(mix_word_29_), .in_30_(mix_word_30_), .in_31_(mix_word_31_), .outx_0_(outx_0_), .outx_1_(outx_1_), .outx_2_(outx_2_), .outx_3_(outx_3_), .outx_4_(outx_4_), .outx_5_(outx_5_), .outx_6_(outx_6_), .outx_7_(outx_7_), .outx_8_(outx_8_), .outx_9_(outx_9_), .outx_10_(outx_10_), .outx_11_(outx_11_), .outx_12_(outx_12_), .outx_13_(outx_13_), .outx_14_(outx_14_), .outx_15_(outx_15_), .outx_16_(outx_16_), .outx_17_(outx_17_), .outx_18_(outx_18_), .outx_19_(outx_19_), .outx_20_(outx_20_), .outx_21_(outx_21_), .outx_22_(outx_22_), .outx_23_(outx_23_), .outx_24_(outx_24_), .outx_25_(outx_25_), .outx_26_(outx_26_), .outx_27_(outx_27_), .outx_28_(outx_28_), .outx_29_(outx_29_), .outx_30_(outx_30_), .outx_31_(outx_31_), .outy_0_(outy_0_), .outy_1_(outy_1_), .outy_2_(outy_2_), .outy_3_(outy_3_), .outy_4_(outy_4_), .outy_5_(outy_5_), .outy_6_(outy_6_), .outy_7_(outy_7_), .outy_8_(outy_8_), .outy_9_(outy_9_), .outy_10_(outy_10_), .outy_11_(outy_11_), .outy_12_(outy_12_), .outy_13_(outy_13_), .outy_14_(outy_14_), .outy_15_(outy_15_), .outy_16_(outy_16_), .outy_17_(outy_17_), .outy_18_(outy_18_), .outy_19_(outy_19_), .outy_20_(outy_20_), .outy_21_(outy_21_), .outy_22_(outy_22_), .outy_23_(outy_23_), .outy_24_(outy_24_), .outy_25_(outy_25_), .outy_26_(outy_26_), .outy_27_(outy_27_), .outy_28_(outy_28_), .outy_29_(outy_29_), .outy_30_(outy_30_), .outy_31_(outy_31_));
endmodule

module word_mixcolum (in_0_, in_1_, in_2_, in_3_, in_4_, in_5_, in_6_, in_7_, in_8_, in_9_, in_10_, in_11_, in_12_, in_13_, in_14_, in_15_, in_16_, in_17_, in_18_, in_19_, in_20_, in_21_, in_22_, in_23_, in_24_, in_25_, in_26_, in_27_, in_28_, in_29_, in_30_, in_31_, outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outx_8_, outx_9_, outx_10_, outx_11_, outx_12_, outx_13_, outx_14_, outx_15_, outx_16_, outx_17_, outx_18_, outx_19_, outx_20_, outx_21_, outx_22_, outx_23_, outx_24_, outx_25_, outx_26_, outx_27_, outx_28_, outx_29_, outx_30_, outx_31_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_, outy_8_, outy_9_, outy_10_, outy_11_, outy_12_, outy_13_, outy_14_, outy_15_, outy_16_, outy_17_, outy_18_, outy_19_, outy_20_, outy_21_, outy_22_, outy_23_, outy_24_, outy_25_, outy_26_, outy_27_, outy_28_, outy_29_, outy_30_, outy_31_);
input in_0_, in_1_, in_2_, in_3_, in_4_, in_5_, in_6_, in_7_, in_8_, in_9_, in_10_, in_11_, in_12_, in_13_, in_14_, in_15_, in_16_, in_17_, in_18_, in_19_, in_20_, in_21_, in_22_, in_23_, in_24_, in_25_, in_26_, in_27_, in_28_, in_29_, in_30_, in_31_;
output outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outx_8_, outx_9_, outx_10_, outx_11_, outx_12_, outx_13_, outx_14_, outx_15_, outx_16_, outx_17_, outx_18_, outx_19_, outx_20_, outx_21_, outx_22_, outx_23_, outx_24_, outx_25_, outx_26_, outx_27_, outx_28_, outx_29_, outx_30_, outx_31_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_, outy_8_, outy_9_, outy_10_, outy_11_, outy_12_, outy_13_, outy_14_, outy_15_, outy_16_, outy_17_, outy_18_, outy_19_, outy_20_, outy_21_, outy_22_, outy_23_, outy_24_, outy_25_, outy_26_, outy_27_, outy_28_, outy_29_, outy_30_, outy_31_;

sg13g2_inv_4 U1 (.A(n14), .Y(n15));
sg13g2_inv_4 U2 (.A(in_23_), .Y(n1));
sg13g2_inv_4 U3 (.A(n1), .Y(n2));
sg13g2_inv_4 U4 (.A(in_13_), .Y(n3));
sg13g2_inv_4 U5 (.A(n3), .Y(n4));
sg13g2_inv_4 U6 (.A(in_15_), .Y(n5));
sg13g2_inv_4 U7 (.A(n5), .Y(n6));
sg13g2_inv_4 U8 (.A(in_29_), .Y(n7));
sg13g2_inv_4 U9 (.A(n7), .Y(n8));
sg13g2_buf_8 U10 (.A(in_24_), .X(n9));
sg13g2_inv_4 U11 (.A(in_7_), .Y(n10));
sg13g2_inv_4 U12 (.A(n10), .Y(n11));
sg13g2_inv_4 U13 (.A(in_31_), .Y(n12));
sg13g2_inv_4 U14 (.A(n12), .Y(n13));
sg13g2_inv_4 U15 (.A(in_21_), .Y(n14));
sg13g2_buf_8 U16 (.A(in_16_), .X(n16));
sg13g2_buf_8 U17 (.A(in_14_), .X(n17));
sg13g2_buf_8 U18 (.A(in_6_), .X(n18));
sg13g2_buf_8 U19 (.A(in_30_), .X(n19));
sg13g2_inv_4 U20 (.A(in_5_), .Y(n20));
sg13g2_inv_4 U21 (.A(n20), .Y(n21));
sg13g2_buf_8 U22 (.A(in_22_), .X(n22));
byte_mixcolum_0 bm1(.a_0_(in_24_), .a_1_(in_25_), .a_2_(in_26_), .a_3_(in_27_), .a_4_(in_28_), .a_5_(n8), .a_6_(n19), .a_7_(n13), .b_0_(n16), .b_1_(in_17_), .b_2_(in_18_), .b_3_(in_19_), .b_4_(in_20_), .b_5_(n15), .b_6_(in_22_), .b_7_(n2), .c_0_(in_8_), .c_1_(in_9_), .c_2_(in_10_), .c_3_(in_11_), .c_4_(in_12_), .c_5_(n4), .c_6_(n17), .c_7_(n6), .d_0_(in_0_), .d_1_(in_1_), .d_2_(in_2_), .d_3_(in_3_), .d_4_(in_4_), .d_5_(n21), .d_6_(n18), .d_7_(n11), .outx_0_(outx_24_), .outx_1_(outx_25_), .outx_2_(outx_26_), .outx_3_(outx_27_), .outx_4_(outx_28_), .outx_5_(outx_29_), .outx_6_(outx_30_), .outx_7_(outx_31_), .outy_0_(outy_24_), .outy_1_(outy_25_), .outy_2_(outy_26_), .outy_3_(outy_27_), .outy_4_(outy_28_), .outy_5_(outy_29_), .outy_6_(outy_30_), .outy_7_(outy_31_));
byte_mixcolum_3 bm2(.a_0_(in_16_), .a_1_(in_17_), .a_2_(in_18_), .a_3_(in_19_), .a_4_(in_20_), .a_5_(n15), .a_6_(n22), .a_7_(n2), .b_0_(in_8_), .b_1_(in_9_), .b_2_(in_10_), .b_3_(in_11_), .b_4_(in_12_), .b_5_(n4), .b_6_(in_14_), .b_7_(n6), .c_0_(in_0_), .c_1_(in_1_), .c_2_(in_2_), .c_3_(in_3_), .c_4_(in_4_), .c_5_(n21), .c_6_(n18), .c_7_(n11), .d_0_(in_24_), .d_1_(in_25_), .d_2_(in_26_), .d_3_(in_27_), .d_4_(in_28_), .d_5_(n8), .d_6_(n19), .d_7_(n13), .outx_0_(outx_16_), .outx_1_(outx_17_), .outx_2_(outx_18_), .outx_3_(outx_19_), .outx_4_(outx_20_), .outx_5_(outx_21_), .outx_6_(outx_22_), .outx_7_(outx_23_), .outy_0_(outy_16_), .outy_1_(outy_17_), .outy_2_(outy_18_), .outy_3_(outy_19_), .outy_4_(outy_20_), .outy_5_(outy_21_), .outy_6_(outy_22_), .outy_7_(outy_23_));
byte_mixcolum_2 bm3(.a_0_(in_8_), .a_1_(in_9_), .a_2_(in_10_), .a_3_(in_11_), .a_4_(in_12_), .a_5_(n4), .a_6_(n17), .a_7_(n6), .b_0_(in_0_), .b_1_(in_1_), .b_2_(in_2_), .b_3_(in_3_), .b_4_(in_4_), .b_5_(n21), .b_6_(in_6_), .b_7_(n11), .c_0_(n9), .c_1_(in_25_), .c_2_(in_26_), .c_3_(in_27_), .c_4_(in_28_), .c_5_(n8), .c_6_(n19), .c_7_(n13), .d_0_(n16), .d_1_(in_17_), .d_2_(in_18_), .d_3_(in_19_), .d_4_(in_20_), .d_5_(n15), .d_6_(n22), .d_7_(n2), .outx_0_(outx_8_), .outx_1_(outx_9_), .outx_2_(outx_10_), .outx_3_(outx_11_), .outx_4_(outx_12_), .outx_5_(outx_13_), .outx_6_(outx_14_), .outx_7_(outx_15_), .outy_0_(outy_8_), .outy_1_(outy_9_), .outy_2_(outy_10_), .outy_3_(outy_11_), .outy_4_(outy_12_), .outy_5_(outy_13_), .outy_6_(outy_14_), .outy_7_(outy_15_));
byte_mixcolum_1 bm4(.a_0_(in_0_), .a_1_(in_1_), .a_2_(in_2_), .a_3_(in_3_), .a_4_(in_4_), .a_5_(n21), .a_6_(in_6_), .a_7_(n11), .b_0_(n9), .b_1_(in_25_), .b_2_(in_26_), .b_3_(in_27_), .b_4_(in_28_), .b_5_(n8), .b_6_(in_30_), .b_7_(n13), .c_0_(n16), .c_1_(in_17_), .c_2_(in_18_), .c_3_(in_19_), .c_4_(in_20_), .c_5_(n15), .c_6_(n22), .c_7_(n2), .d_0_(in_8_), .d_1_(in_9_), .d_2_(in_10_), .d_3_(in_11_), .d_4_(in_12_), .d_5_(n4), .d_6_(n17), .d_7_(n6), .outx_0_(outx_0_), .outx_1_(outx_1_), .outx_2_(outx_2_), .outx_3_(outx_3_), .outx_4_(outx_4_), .outx_5_(outx_5_), .outx_6_(outx_6_), .outx_7_(outx_7_), .outy_0_(outy_0_), .outy_1_(outy_1_), .outy_2_(outy_2_), .outy_3_(outy_3_), .outy_4_(outy_4_), .outy_5_(outy_5_), .outy_6_(outy_6_), .outy_7_(outy_7_));
endmodule

module byte_mixcolum_1 (a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_);
input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
output outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_;

sg13g2_inv_4 U1 (.A(n146), .Y(outy_7_));
sg13g2_xnor2_1 U2 (.A(n145), .B(n144), .Y(n146));
sg13g2_xnor2_1 U3 (.A(n143), .B(n142), .Y(n144));
sg13g2_xnor2_1 U4 (.A(n141), .B(n140), .Y(n142));
sg13g2_xnor2_1 U5 (.A(c_4_), .B(n139), .Y(n145));
sg13g2_xnor2_1 U6 (.A(d_4_), .B(c_5_), .Y(n139));
sg13g2_xnor2_1 U7 (.A(n138), .B(n137), .Y(outy_6_));
sg13g2_xnor2_1 U8 (.A(n136), .B(n135), .Y(n137));
sg13g2_xnor2_1 U9 (.A(n134), .B(n133), .Y(n136));
sg13g2_xnor2_1 U10 (.A(a_4_), .B(n132), .Y(n138));
sg13g2_xnor2_1 U11 (.A(d_7_), .B(a_7_), .Y(n132));
sg13g2_xnor2_1 U12 (.A(n131), .B(n130), .Y(outy_5_));
sg13g2_xnor2_1 U13 (.A(n129), .B(n128), .Y(n130));
sg13g2_xnor2_1 U14 (.A(n143), .B(n127), .Y(n129));
sg13g2_xnor2_1 U15 (.A(n126), .B(n125), .Y(n131));
sg13g2_xnor2_1 U16 (.A(c_2_), .B(a_3_), .Y(n125));
sg13g2_xnor2_1 U17 (.A(d_2_), .B(c_3_), .Y(n126));
sg13g2_xnor2_1 U18 (.A(n124), .B(n123), .Y(outy_4_));
sg13g2_xnor2_1 U19 (.A(n122), .B(n135), .Y(n123));
sg13g2_xnor2_1 U20 (.A(b_1_), .B(n103), .Y(n98));
sg13g2_xnor2_1 U21 (.A(c_1_), .B(a_2_), .Y(n122));
sg13g2_xnor2_1 U22 (.A(n119), .B(n118), .Y(n124));
sg13g2_xnor2_1 U23 (.A(n117), .B(n116), .Y(n118));
sg13g2_xnor2_1 U24 (.A(b_1_), .B(n96), .Y(n117));
sg13g2_xnor2_1 U25 (.A(c_6_), .B(n91), .Y(n109));
sg13g2_xnor2_1 U26 (.A(d_1_), .B(n91), .Y(n116));
sg13g2_xnor2_1 U27 (.A(n121), .B(n120), .Y(n135));
sg13g2_inv_4 U28 (.A(n108), .Y(n110));
sg13g2_xnor2_1 U29 (.A(c_4_), .B(a_3_), .Y(n121));
sg13g2_xnor2_1 U30 (.A(n141), .B(n134), .Y(n106));
sg13g2_xnor2_1 U31 (.A(n105), .B(n104), .Y(n141));
sg13g2_xnor2_1 U32 (.A(a_1_), .B(n103), .Y(n107));
sg13g2_xnor2_1 U33 (.A(n102), .B(n101), .Y(outy_2_));
sg13g2_xnor2_1 U34 (.A(n100), .B(n127), .Y(n101));
sg13g2_xnor2_1 U35 (.A(c_7_), .B(a_5_), .Y(n104));
sg13g2_xnor2_1 U36 (.A(c_6_), .B(c_0_), .Y(n100));
sg13g2_xnor2_1 U37 (.A(n98), .B(n97), .Y(n102));
sg13g2_xnor2_1 U38 (.A(n96), .B(n95), .Y(n97));
sg13g2_xnor2_1 U39 (.A(n94), .B(n93), .Y(outy_1_));
sg13g2_xnor2_1 U40 (.A(n116), .B(n120), .Y(n93));
sg13g2_xnor2_1 U41 (.A(c_2_), .B(a_1_), .Y(n96));
sg13g2_xnor2_1 U42 (.A(b_0_), .B(n111), .Y(n74));
sg13g2_inv_4 U43 (.A(n104), .Y(n92));
sg13g2_xnor2_1 U44 (.A(d_3_), .B(c_3_), .Y(n77));
sg13g2_xnor2_1 U45 (.A(n107), .B(n106), .Y(n115));
sg13g2_xnor2_1 U46 (.A(n90), .B(n89), .Y(outy_0_));
sg13g2_xnor2_1 U47 (.A(n109), .B(outx_0_), .Y(n89));
sg13g2_xnor2_1 U48 (.A(b_7_), .B(a_7_), .Y(n81));
sg13g2_xnor2_1 U49 (.A(a_6_), .B(a_5_), .Y(n90));
sg13g2_xnor2_1 U50 (.A(n88), .B(n140), .Y(outx_7_));
sg13g2_inv_4 U51 (.A(a_0_), .Y(n103));
sg13g2_xnor2_1 U52 (.A(n86), .B(n105), .Y(n88));
sg13g2_xnor2_1 U53 (.A(n81), .B(n74), .Y(outx_0_));
sg13g2_inv_4 U54 (.A(c_7_), .Y(n86));
sg13g2_xnor2_1 U55 (.A(n85), .B(n84), .Y(outx_6_));
sg13g2_xnor2_1 U56 (.A(n87), .B(d_6_), .Y(n84));
sg13g2_xnor2_1 U57 (.A(d_0_), .B(c_0_), .Y(n111));
sg13g2_xnor2_1 U58 (.A(n83), .B(n133), .Y(n85));
sg13g2_xnor2_1 U59 (.A(c_6_), .B(b_5_), .Y(n133));
sg13g2_inv_4 U60 (.A(a_5_), .Y(n83));
sg13g2_xnor2_1 U61 (.A(n143), .B(n91), .Y(outx_5_));
sg13g2_xnor2_1 U62 (.A(c_5_), .B(d_5_), .Y(n82));
sg13g2_xnor2_1 U63 (.A(c_1_), .B(b_0_), .Y(n113));
sg13g2_xnor2_1 U64 (.A(b_4_), .B(a_4_), .Y(n143));
sg13g2_xnor2_1 U65 (.A(n81), .B(n80), .Y(outx_4_));
sg13g2_xnor2_1 U66 (.A(n121), .B(n119), .Y(n80));
sg13g2_xnor2_1 U67 (.A(b_3_), .B(n79), .Y(n119));
sg13g2_xnor2_1 U68 (.A(d_4_), .B(b_4_), .Y(n79));
sg13g2_xnor2_1 U69 (.A(n115), .B(n114), .Y(outy_3_));
sg13g2_xnor2_1 U70 (.A(n81), .B(n78), .Y(outx_3_));
sg13g2_xnor2_1 U71 (.A(n108), .B(n134), .Y(n78));
sg13g2_xnor2_1 U72 (.A(n105), .B(n99), .Y(n127));
sg13g2_xnor2_1 U73 (.A(b_3_), .B(n77), .Y(n134));
sg13g2_xnor2_1 U74 (.A(b_2_), .B(a_2_), .Y(n108));
sg13g2_xnor2_1 U75 (.A(n95), .B(n117), .Y(outx_2_));
sg13g2_xnor2_1 U76 (.A(n113), .B(n112), .Y(n114));
sg13g2_xnor2_1 U77 (.A(d_7_), .B(a_6_), .Y(n105));
sg13g2_xnor2_1 U78 (.A(d_2_), .B(b_2_), .Y(n95));
sg13g2_xnor2_1 U79 (.A(n76), .B(n81), .Y(outx_1_));
sg13g2_xnor2_1 U80 (.A(d_1_), .B(n94), .Y(n76));
sg13g2_inv_4 U81 (.A(n75), .Y(n94));
sg13g2_xnor2_1 U82 (.A(n113), .B(n98), .Y(n75));
sg13g2_xnor2_1 U83 (.A(n111), .B(n128), .Y(n112));
sg13g2_xnor2_1 U84 (.A(d_6_), .B(n140), .Y(n99));
sg13g2_inv_4 U85 (.A(b_6_), .Y(n87));
sg13g2_xnor2_1 U86 (.A(n92), .B(n99), .Y(n120));
sg13g2_xnor2_1 U87 (.A(b_5_), .B(n82), .Y(n91));
sg13g2_xnor2_1 U88 (.A(n110), .B(n109), .Y(n128));
sg13g2_xnor2_1 U89 (.A(n87), .B(b_7_), .Y(n140));
endmodule

module byte_mixcolum_3 (a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_);
input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
output outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_;

sg13g2_xnor2_1 U1 (.A(n117), .B(n118), .Y(n119));
sg13g2_xnor2_1 U2 (.A(n145), .B(n146), .Y(n147));
sg13g2_xnor2_1 U3 (.A(n143), .B(n144), .Y(n145));
sg13g2_xnor2_1 U4 (.A(n142), .B(n141), .Y(n143));
sg13g2_xnor2_1 U5 (.A(c_4_), .B(n140), .Y(n146));
sg13g2_xnor2_1 U6 (.A(d_4_), .B(c_5_), .Y(n140));
sg13g2_xnor2_1 U7 (.A(b_1_), .B(n97), .Y(n118));
sg13g2_xnor2_1 U8 (.A(n114), .B(n99), .Y(n76));
sg13g2_xnor2_1 U9 (.A(n135), .B(n134), .Y(n137));
sg13g2_xnor2_1 U10 (.A(a_4_), .B(n133), .Y(n139));
sg13g2_xnor2_1 U11 (.A(d_7_), .B(a_7_), .Y(n133));
sg13g2_xnor2_1 U12 (.A(b_1_), .B(n104), .Y(n99));
sg13g2_xnor2_1 U13 (.A(n123), .B(n136), .Y(n124));
sg13g2_xnor2_1 U14 (.A(n139), .B(n138), .Y(outy_6_));
sg13g2_xnor2_1 U15 (.A(n127), .B(n126), .Y(n132));
sg13g2_xnor2_1 U16 (.A(c_2_), .B(a_3_), .Y(n126));
sg13g2_xnor2_1 U17 (.A(d_2_), .B(c_3_), .Y(n127));
sg13g2_xnor2_1 U18 (.A(n125), .B(n124), .Y(outy_4_));
sg13g2_xnor2_1 U19 (.A(n137), .B(n136), .Y(n138));
sg13g2_xnor2_1 U20 (.A(n116), .B(n115), .Y(outy_3_));
sg13g2_xnor2_1 U21 (.A(c_1_), .B(a_2_), .Y(n123));
sg13g2_xnor2_1 U22 (.A(n119), .B(n120), .Y(n125));
sg13g2_xnor2_1 U23 (.A(b_4_), .B(a_4_), .Y(n144));
sg13g2_xnor2_1 U24 (.A(n106), .B(n100), .Y(n128));
sg13g2_xnor2_1 U25 (.A(b_7_), .B(n88), .Y(n141));
sg13g2_xnor2_1 U26 (.A(n132), .B(n131), .Y(outy_5_));
sg13g2_xnor2_1 U27 (.A(n130), .B(n129), .Y(n131));
sg13g2_inv_4 U28 (.A(n109), .Y(n111));
sg13g2_xnor2_1 U29 (.A(n108), .B(n107), .Y(n116));
sg13g2_xnor2_1 U30 (.A(n142), .B(n135), .Y(n107));
sg13g2_xnor2_1 U31 (.A(n105), .B(n106), .Y(n142));
sg13g2_xnor2_1 U32 (.A(a_1_), .B(n104), .Y(n108));
sg13g2_xnor2_1 U33 (.A(n103), .B(n102), .Y(outy_2_));
sg13g2_xnor2_1 U34 (.A(n101), .B(n128), .Y(n102));
sg13g2_xnor2_1 U35 (.A(n111), .B(n110), .Y(n129));
sg13g2_xnor2_1 U36 (.A(c_6_), .B(c_0_), .Y(n101));
sg13g2_xnor2_1 U37 (.A(n99), .B(n98), .Y(n103));
sg13g2_xnor2_1 U38 (.A(n97), .B(n96), .Y(n98));
sg13g2_xnor2_1 U39 (.A(n95), .B(n94), .Y(outy_1_));
sg13g2_xnor2_1 U40 (.A(n117), .B(n121), .Y(n94));
sg13g2_xnor2_1 U41 (.A(n144), .B(n128), .Y(n130));
sg13g2_xnor2_1 U42 (.A(c_2_), .B(a_1_), .Y(n97));
sg13g2_inv_4 U43 (.A(n105), .Y(n93));
sg13g2_xnor2_1 U44 (.A(c_7_), .B(a_5_), .Y(n105));
sg13g2_inv_4 U45 (.A(n147), .Y(outy_7_));
sg13g2_xnor2_1 U46 (.A(n91), .B(n90), .Y(outy_0_));
sg13g2_xnor2_1 U47 (.A(n110), .B(outx_0_), .Y(n90));
sg13g2_xnor2_1 U48 (.A(n74), .B(n75), .Y(outx_0_));
sg13g2_xnor2_1 U49 (.A(a_6_), .B(a_5_), .Y(n91));
sg13g2_xnor2_1 U50 (.A(n89), .B(n141), .Y(outx_7_));
sg13g2_xnor2_1 U51 (.A(b_0_), .B(n112), .Y(n75));
sg13g2_xnor2_1 U52 (.A(n106), .B(n87), .Y(n89));
sg13g2_xnor2_1 U53 (.A(d_1_), .B(n92), .Y(n117));
sg13g2_inv_4 U54 (.A(c_7_), .Y(n87));
sg13g2_xnor2_1 U55 (.A(n86), .B(n85), .Y(outx_6_));
sg13g2_xnor2_1 U56 (.A(n88), .B(d_6_), .Y(n85));
sg13g2_xnor2_1 U57 (.A(c_1_), .B(b_0_), .Y(n114));
sg13g2_xnor2_1 U58 (.A(n84), .B(n134), .Y(n86));
sg13g2_xnor2_1 U59 (.A(c_6_), .B(b_5_), .Y(n134));
sg13g2_inv_4 U60 (.A(a_5_), .Y(n84));
sg13g2_xnor2_1 U61 (.A(n144), .B(n92), .Y(outx_5_));
sg13g2_xnor2_1 U62 (.A(b_5_), .B(n83), .Y(n92));
sg13g2_xnor2_1 U63 (.A(d_7_), .B(a_6_), .Y(n106));
sg13g2_xnor2_1 U64 (.A(d_0_), .B(c_0_), .Y(n112));
sg13g2_xnor2_1 U65 (.A(n74), .B(n81), .Y(outx_4_));
sg13g2_xnor2_1 U66 (.A(n122), .B(n120), .Y(n81));
sg13g2_xnor2_1 U67 (.A(b_3_), .B(n80), .Y(n120));
sg13g2_xnor2_1 U68 (.A(d_4_), .B(b_4_), .Y(n80));
sg13g2_xnor2_1 U69 (.A(n93), .B(n100), .Y(n121));
sg13g2_xnor2_1 U70 (.A(n74), .B(n79), .Y(outx_3_));
sg13g2_xnor2_1 U71 (.A(n109), .B(n135), .Y(n79));
sg13g2_xnor2_1 U72 (.A(d_6_), .B(n141), .Y(n100));
sg13g2_xnor2_1 U73 (.A(n114), .B(n113), .Y(n115));
sg13g2_xnor2_1 U74 (.A(b_2_), .B(a_2_), .Y(n109));
sg13g2_xnor2_1 U75 (.A(n96), .B(n118), .Y(outx_2_));
sg13g2_buf_8 U76 (.A(n82), .X(n74));
sg13g2_xnor2_1 U77 (.A(n112), .B(n129), .Y(n113));
sg13g2_xnor2_1 U78 (.A(d_2_), .B(b_2_), .Y(n96));
sg13g2_xnor2_1 U79 (.A(n77), .B(n74), .Y(outx_1_));
sg13g2_xnor2_1 U80 (.A(d_1_), .B(n95), .Y(n77));
sg13g2_inv_4 U81 (.A(n76), .Y(n95));
sg13g2_xnor2_1 U82 (.A(c_4_), .B(a_3_), .Y(n122));
sg13g2_inv_4 U83 (.A(b_6_), .Y(n88));
sg13g2_inv_4 U84 (.A(a_0_), .Y(n104));
sg13g2_xnor2_1 U85 (.A(d_5_), .B(c_5_), .Y(n83));
sg13g2_xnor2_1 U86 (.A(d_3_), .B(c_3_), .Y(n78));
sg13g2_xnor2_1 U87 (.A(b_3_), .B(n78), .Y(n135));
sg13g2_xnor2_1 U88 (.A(c_6_), .B(n92), .Y(n110));
sg13g2_xnor2_1 U89 (.A(b_7_), .B(a_7_), .Y(n82));
sg13g2_xnor2_1 U90 (.A(n122), .B(n121), .Y(n136));
endmodule

module byte_mixcolum_2 (a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_);
input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
output outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_;

sg13g2_inv_4 U1 (.A(n147), .Y(outy_7_));
sg13g2_xnor2_1 U2 (.A(n146), .B(n145), .Y(n147));
sg13g2_xnor2_1 U3 (.A(n144), .B(n74), .Y(outx_5_));
sg13g2_xnor2_1 U4 (.A(n144), .B(n143), .Y(n145));
sg13g2_xnor2_1 U5 (.A(c_4_), .B(n140), .Y(n146));
sg13g2_xnor2_1 U6 (.A(c_5_), .B(d_4_), .Y(n140));
sg13g2_xnor2_1 U7 (.A(b_4_), .B(a_4_), .Y(n144));
sg13g2_xnor2_1 U8 (.A(b_7_), .B(n88), .Y(n141));
sg13g2_inv_4 U9 (.A(b_6_), .Y(n88));
sg13g2_xnor2_1 U10 (.A(a_4_), .B(n133), .Y(n139));
sg13g2_xnor2_1 U11 (.A(d_7_), .B(a_7_), .Y(n133));
sg13g2_xnor2_1 U12 (.A(n132), .B(n131), .Y(outy_5_));
sg13g2_xnor2_1 U13 (.A(n130), .B(n129), .Y(n131));
sg13g2_xnor2_1 U14 (.A(n93), .B(n100), .Y(n121));
sg13g2_xnor2_1 U15 (.A(n127), .B(n126), .Y(n132));
sg13g2_xnor2_1 U16 (.A(c_2_), .B(a_3_), .Y(n126));
sg13g2_xnor2_1 U17 (.A(d_2_), .B(c_3_), .Y(n127));
sg13g2_xnor2_1 U18 (.A(n144), .B(n128), .Y(n130));
sg13g2_xnor2_1 U19 (.A(b_1_), .B(n97), .Y(n118));
sg13g2_buf_8 U20 (.A(n92), .X(n74));
sg13g2_xnor2_1 U21 (.A(c_1_), .B(a_2_), .Y(n123));
sg13g2_xnor2_1 U22 (.A(n119), .B(n120), .Y(n125));
sg13g2_xnor2_1 U23 (.A(n118), .B(n117), .Y(n119));
sg13g2_xnor2_1 U24 (.A(n123), .B(n136), .Y(n124));
sg13g2_xnor2_1 U25 (.A(n114), .B(n113), .Y(n115));
sg13g2_xnor2_1 U26 (.A(n135), .B(n134), .Y(n137));
sg13g2_xnor2_1 U27 (.A(n142), .B(n141), .Y(n143));
sg13g2_xnor2_1 U28 (.A(c_2_), .B(a_1_), .Y(n97));
sg13g2_xnor2_1 U29 (.A(n108), .B(n107), .Y(n116));
sg13g2_xnor2_1 U30 (.A(n142), .B(n135), .Y(n107));
sg13g2_xnor2_1 U31 (.A(d_0_), .B(c_0_), .Y(n112));
sg13g2_xnor2_1 U32 (.A(n104), .B(a_1_), .Y(n108));
sg13g2_xnor2_1 U33 (.A(n103), .B(n102), .Y(outy_2_));
sg13g2_xnor2_1 U34 (.A(n101), .B(n128), .Y(n102));
sg13g2_xnor2_1 U35 (.A(n112), .B(n129), .Y(n113));
sg13g2_xnor2_1 U36 (.A(c_6_), .B(c_0_), .Y(n101));
sg13g2_xnor2_1 U37 (.A(n99), .B(n98), .Y(n103));
sg13g2_xnor2_1 U38 (.A(n97), .B(n96), .Y(n98));
sg13g2_xnor2_1 U39 (.A(n95), .B(n94), .Y(outy_1_));
sg13g2_xnor2_1 U40 (.A(n117), .B(n121), .Y(n94));
sg13g2_xnor2_1 U41 (.A(n106), .B(n105), .Y(n142));
sg13g2_inv_4 U42 (.A(n105), .Y(n93));
sg13g2_xnor2_1 U43 (.A(c_7_), .B(a_5_), .Y(n105));
sg13g2_xnor2_1 U44 (.A(b_7_), .B(a_7_), .Y(n82));
sg13g2_xnor2_1 U45 (.A(b_1_), .B(n104), .Y(n99));
sg13g2_xnor2_1 U46 (.A(n91), .B(n90), .Y(outy_0_));
sg13g2_xnor2_1 U47 (.A(n110), .B(outx_0_), .Y(n90));
sg13g2_inv_4 U48 (.A(a_0_), .Y(n104));
sg13g2_xnor2_1 U49 (.A(a_6_), .B(a_5_), .Y(n91));
sg13g2_xnor2_1 U50 (.A(n89), .B(n141), .Y(outx_7_));
sg13g2_xnor2_1 U51 (.A(d_1_), .B(n92), .Y(n117));
sg13g2_xnor2_1 U52 (.A(n87), .B(n106), .Y(n89));
sg13g2_xnor2_1 U53 (.A(n125), .B(n124), .Y(outy_4_));
sg13g2_inv_4 U54 (.A(c_7_), .Y(n87));
sg13g2_xnor2_1 U55 (.A(n86), .B(n85), .Y(outx_6_));
sg13g2_xnor2_1 U56 (.A(n88), .B(d_6_), .Y(n85));
sg13g2_xnor2_1 U57 (.A(n115), .B(n116), .Y(outy_3_));
sg13g2_xnor2_1 U58 (.A(n84), .B(n134), .Y(n86));
sg13g2_xnor2_1 U59 (.A(c_6_), .B(b_5_), .Y(n134));
sg13g2_inv_4 U60 (.A(a_5_), .Y(n84));
sg13g2_xnor2_1 U61 (.A(n106), .B(n100), .Y(n128));
sg13g2_xnor2_1 U62 (.A(d_6_), .B(n141), .Y(n100));
sg13g2_xnor2_1 U63 (.A(n111), .B(n110), .Y(n129));
sg13g2_xnor2_1 U64 (.A(n139), .B(n138), .Y(outy_6_));
sg13g2_xnor2_1 U65 (.A(n82), .B(n81), .Y(outx_4_));
sg13g2_xnor2_1 U66 (.A(n122), .B(n120), .Y(n81));
sg13g2_xnor2_1 U67 (.A(n137), .B(n136), .Y(n138));
sg13g2_xnor2_1 U68 (.A(b_5_), .B(n83), .Y(n92));
sg13g2_xnor2_1 U69 (.A(c_4_), .B(a_3_), .Y(n122));
sg13g2_xnor2_1 U70 (.A(n82), .B(n79), .Y(outx_3_));
sg13g2_xnor2_1 U71 (.A(n109), .B(n135), .Y(n79));
sg13g2_xnor2_1 U72 (.A(d_4_), .B(b_4_), .Y(n80));
sg13g2_xnor2_1 U73 (.A(b_3_), .B(n80), .Y(n120));
sg13g2_xnor2_1 U74 (.A(d_5_), .B(c_5_), .Y(n83));
sg13g2_xnor2_1 U75 (.A(n96), .B(n118), .Y(outx_2_));
sg13g2_xnor2_1 U76 (.A(b_0_), .B(n112), .Y(n75));
sg13g2_inv_4 U77 (.A(n109), .Y(n111));
sg13g2_xnor2_1 U78 (.A(d_2_), .B(b_2_), .Y(n96));
sg13g2_xnor2_1 U79 (.A(n77), .B(n82), .Y(outx_1_));
sg13g2_xnor2_1 U80 (.A(d_1_), .B(n95), .Y(n77));
sg13g2_inv_4 U81 (.A(n76), .Y(n95));
sg13g2_xnor2_1 U82 (.A(n114), .B(n99), .Y(n76));
sg13g2_xnor2_1 U83 (.A(b_2_), .B(a_2_), .Y(n109));
sg13g2_xnor2_1 U84 (.A(b_3_), .B(n78), .Y(n135));
sg13g2_xnor2_1 U85 (.A(c_1_), .B(b_0_), .Y(n114));
sg13g2_xnor2_1 U86 (.A(d_3_), .B(c_3_), .Y(n78));
sg13g2_xnor2_1 U87 (.A(n92), .B(c_6_), .Y(n110));
sg13g2_xnor2_1 U88 (.A(n82), .B(n75), .Y(outx_0_));
sg13g2_xnor2_1 U89 (.A(d_7_), .B(a_6_), .Y(n106));
sg13g2_xnor2_1 U90 (.A(n122), .B(n121), .Y(n136));
endmodule

module byte_mixcolum_0 (a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_);
input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
output outx_0_, outx_1_, outx_2_, outx_3_, outx_4_, outx_5_, outx_6_, outx_7_, outy_0_, outy_1_, outy_2_, outy_3_, outy_4_, outy_5_, outy_6_, outy_7_;

sg13g2_xnor2_1 U1 (.A(n40), .B(n41), .Y(n32));
sg13g2_xnor2_1 U2 (.A(n3), .B(n2), .Y(n1));
sg13g2_xnor2_1 U3 (.A(n4), .B(n5), .Y(n3));
sg13g2_xnor2_1 U4 (.A(n6), .B(n7), .Y(n5));
sg13g2_xnor2_1 U5 (.A(c_4_), .B(n8), .Y(n2));
sg13g2_xnor2_1 U6 (.A(d_4_), .B(c_5_), .Y(n8));
sg13g2_xnor2_1 U7 (.A(n4), .B(n20), .Y(n18));
sg13g2_inv_4 U8 (.A(c_7_), .Y(n61));
sg13g2_xnor2_1 U9 (.A(n13), .B(n14), .Y(n11));
sg13g2_xnor2_1 U10 (.A(a_4_), .B(n15), .Y(n9));
sg13g2_xnor2_1 U11 (.A(d_7_), .B(a_7_), .Y(n15));
sg13g2_xnor2_1 U12 (.A(n17), .B(n16), .Y(outy_5_));
sg13g2_xnor2_1 U13 (.A(n18), .B(n19), .Y(n17));
sg13g2_xnor2_1 U14 (.A(b_5_), .B(n65), .Y(n56));
sg13g2_xnor2_1 U15 (.A(n21), .B(n22), .Y(n16));
sg13g2_xnor2_1 U16 (.A(c_2_), .B(a_3_), .Y(n22));
sg13g2_xnor2_1 U17 (.A(d_2_), .B(c_3_), .Y(n21));
sg13g2_xnor2_1 U18 (.A(d_5_), .B(c_5_), .Y(n65));
sg13g2_xnor2_1 U19 (.A(n42), .B(n43), .Y(n6));
sg13g2_xnor2_1 U20 (.A(d_7_), .B(a_6_), .Y(n42));
sg13g2_xnor2_1 U21 (.A(c_1_), .B(a_2_), .Y(n25));
sg13g2_xnor2_1 U22 (.A(n28), .B(n29), .Y(n23));
sg13g2_xnor2_1 U23 (.A(n37), .B(n38), .Y(n19));
sg13g2_xnor2_1 U24 (.A(c_1_), .B(b_0_), .Y(n34));
sg13g2_xnor2_1 U25 (.A(n30), .B(n31), .Y(n29));
sg13g2_xnor2_1 U26 (.A(b_7_), .B(n60), .Y(n7));
sg13g2_xnor2_1 U27 (.A(n55), .B(n48), .Y(n27));
sg13g2_inv_4 U28 (.A(n39), .Y(n37));
sg13g2_xnor2_1 U29 (.A(n9), .B(n10), .Y(outy_6_));
sg13g2_xnor2_1 U30 (.A(n6), .B(n13), .Y(n41));
sg13g2_xnor2_1 U31 (.A(n11), .B(n12), .Y(n10));
sg13g2_xnor2_1 U32 (.A(n44), .B(a_1_), .Y(n40));
sg13g2_xnor2_1 U33 (.A(n45), .B(n46), .Y(outy_2_));
sg13g2_xnor2_1 U34 (.A(n47), .B(n20), .Y(n46));
sg13g2_xnor2_1 U35 (.A(b_7_), .B(a_7_), .Y(n66));
sg13g2_xnor2_1 U36 (.A(c_6_), .B(c_0_), .Y(n47));
sg13g2_xnor2_1 U37 (.A(n49), .B(n50), .Y(n45));
sg13g2_xnor2_1 U38 (.A(n51), .B(n52), .Y(n50));
sg13g2_xnor2_1 U39 (.A(n54), .B(n53), .Y(outy_1_));
sg13g2_xnor2_1 U40 (.A(n31), .B(n27), .Y(n54));
sg13g2_inv_4 U41 (.A(n1), .Y(outy_7_));
sg13g2_xnor2_1 U42 (.A(d_6_), .B(n7), .Y(n48));
sg13g2_inv_4 U43 (.A(n43), .Y(n55));
sg13g2_xnor2_1 U44 (.A(n24), .B(n23), .Y(outy_4_));
sg13g2_xnor2_1 U45 (.A(n25), .B(n12), .Y(n24));
sg13g2_xnor2_1 U46 (.A(n57), .B(n58), .Y(outy_0_));
sg13g2_xnor2_1 U47 (.A(n38), .B(outx_0_), .Y(n58));
sg13g2_xnor2_1 U48 (.A(n61), .B(n64), .Y(n43));
sg13g2_xnor2_1 U49 (.A(a_6_), .B(a_5_), .Y(n57));
sg13g2_xnor2_1 U50 (.A(n59), .B(n7), .Y(outx_7_));
sg13g2_inv_4 U51 (.A(a_5_), .Y(n64));
sg13g2_xnor2_1 U52 (.A(n61), .B(n42), .Y(n59));
sg13g2_xnor2_1 U53 (.A(b_3_), .B(n70), .Y(n13));
sg13g2_xnor2_1 U54 (.A(d_3_), .B(c_3_), .Y(n70));
sg13g2_xnor2_1 U55 (.A(n62), .B(n63), .Y(outx_6_));
sg13g2_xnor2_1 U56 (.A(n60), .B(d_6_), .Y(n63));
sg13g2_inv_4 U57 (.A(b_6_), .Y(n60));
sg13g2_xnor2_1 U58 (.A(n64), .B(n14), .Y(n62));
sg13g2_xnor2_1 U59 (.A(c_6_), .B(b_5_), .Y(n14));
sg13g2_xnor2_1 U60 (.A(n42), .B(n48), .Y(n20));
sg13g2_xnor2_1 U61 (.A(n4), .B(n56), .Y(outx_5_));
sg13g2_xnor2_1 U62 (.A(d_1_), .B(n56), .Y(n31));
sg13g2_xnor2_1 U63 (.A(b_1_), .B(n51), .Y(n30));
sg13g2_xnor2_1 U64 (.A(b_4_), .B(a_4_), .Y(n4));
sg13g2_xnor2_1 U65 (.A(n66), .B(n67), .Y(outx_4_));
sg13g2_xnor2_1 U66 (.A(n26), .B(n28), .Y(n67));
sg13g2_xnor2_1 U67 (.A(b_3_), .B(n68), .Y(n28));
sg13g2_xnor2_1 U68 (.A(d_4_), .B(b_4_), .Y(n68));
sg13g2_xnor2_1 U69 (.A(c_4_), .B(a_3_), .Y(n26));
sg13g2_xnor2_1 U70 (.A(n66), .B(n69), .Y(outx_3_));
sg13g2_xnor2_1 U71 (.A(n39), .B(n13), .Y(n69));
sg13g2_xnor2_1 U72 (.A(c_2_), .B(a_1_), .Y(n51));
sg13g2_xnor2_1 U73 (.A(n32), .B(n33), .Y(outy_3_));
sg13g2_xnor2_1 U74 (.A(b_2_), .B(a_2_), .Y(n39));
sg13g2_xnor2_1 U75 (.A(n52), .B(n30), .Y(outx_2_));
sg13g2_xnor2_1 U76 (.A(n34), .B(n35), .Y(n33));
sg13g2_xnor2_1 U77 (.A(n66), .B(n73), .Y(outx_0_));
sg13g2_xnor2_1 U78 (.A(d_2_), .B(b_2_), .Y(n52));
sg13g2_xnor2_1 U79 (.A(n71), .B(n66), .Y(outx_1_));
sg13g2_xnor2_1 U80 (.A(d_1_), .B(n53), .Y(n71));
sg13g2_inv_4 U81 (.A(n72), .Y(n53));
sg13g2_xnor2_1 U82 (.A(n49), .B(n34), .Y(n72));
sg13g2_xnor2_1 U83 (.A(b_1_), .B(n44), .Y(n49));
sg13g2_inv_4 U84 (.A(a_0_), .Y(n44));
sg13g2_xnor2_1 U85 (.A(b_0_), .B(n36), .Y(n73));
sg13g2_xnor2_1 U86 (.A(d_0_), .B(c_0_), .Y(n36));
sg13g2_xnor2_1 U87 (.A(n36), .B(n19), .Y(n35));
sg13g2_xnor2_1 U88 (.A(c_6_), .B(n56), .Y(n38));
sg13g2_xnor2_1 U89 (.A(n26), .B(n27), .Y(n12));
endmodule

module keysched192 (clk, last_key_i_0_, last_key_i_1_, last_key_i_2_, last_key_i_3_, last_key_i_4_, last_key_i_5_, last_key_i_6_, last_key_i_7_, last_key_i_8_, last_key_i_9_, last_key_i_10_, last_key_i_11_, last_key_i_12_, last_key_i_13_, last_key_i_14_, last_key_i_15_, last_key_i_16_, last_key_i_17_, last_key_i_18_, last_key_i_19_, last_key_i_20_, last_key_i_21_, last_key_i_22_, last_key_i_23_, last_key_i_24_, last_key_i_25_, last_key_i_26_, last_key_i_27_, last_key_i_28_, last_key_i_29_, last_key_i_30_, last_key_i_31_, last_key_i_32_, last_key_i_33_, last_key_i_34_, last_key_i_35_, last_key_i_36_, last_key_i_37_, last_key_i_38_, last_key_i_39_, last_key_i_40_, last_key_i_41_, last_key_i_42_, last_key_i_43_, last_key_i_44_, last_key_i_45_, last_key_i_46_, last_key_i_47_, last_key_i_48_, last_key_i_49_, last_key_i_50_, last_key_i_51_, last_key_i_52_, last_key_i_53_, last_key_i_54_, last_key_i_55_, last_key_i_56_, last_key_i_57_, last_key_i_58_, last_key_i_59_, last_key_i_60_, last_key_i_61_, last_key_i_62_, last_key_i_63_, last_key_i_64_, last_key_i_65_, last_key_i_66_, last_key_i_67_, last_key_i_68_, last_key_i_69_, last_key_i_70_, last_key_i_71_, last_key_i_72_, last_key_i_73_, last_key_i_74_, last_key_i_75_, last_key_i_76_, last_key_i_77_, last_key_i_78_, last_key_i_79_, last_key_i_80_, last_key_i_81_, last_key_i_82_, last_key_i_83_, last_key_i_84_, last_key_i_85_, last_key_i_86_, last_key_i_87_, last_key_i_88_, last_key_i_89_, last_key_i_90_, last_key_i_91_, last_key_i_92_, last_key_i_93_, last_key_i_94_, last_key_i_95_, last_key_i_96_, last_key_i_97_, last_key_i_98_, last_key_i_99_, last_key_i_100_, last_key_i_101_, last_key_i_102_, last_key_i_103_, last_key_i_104_, last_key_i_105_, last_key_i_106_, last_key_i_107_, last_key_i_108_, last_key_i_109_, last_key_i_110_, last_key_i_111_, last_key_i_112_, last_key_i_113_, last_key_i_114_, last_key_i_115_, last_key_i_116_, last_key_i_117_, last_key_i_118_, last_key_i_119_, last_key_i_120_, last_key_i_121_, last_key_i_122_, last_key_i_123_, last_key_i_124_, last_key_i_125_, last_key_i_126_, last_key_i_127_, last_key_i_128_, last_key_i_129_, last_key_i_130_, last_key_i_131_, last_key_i_132_, last_key_i_133_, last_key_i_134_, last_key_i_135_, last_key_i_136_, last_key_i_137_, last_key_i_138_, last_key_i_139_, last_key_i_140_, last_key_i_141_, last_key_i_142_, last_key_i_143_, last_key_i_144_, last_key_i_145_, last_key_i_146_, last_key_i_147_, last_key_i_148_, last_key_i_149_, last_key_i_150_, last_key_i_151_, last_key_i_152_, last_key_i_153_, last_key_i_154_, last_key_i_155_, last_key_i_156_, last_key_i_157_, last_key_i_158_, last_key_i_159_, last_key_i_160_, last_key_i_161_, last_key_i_162_, last_key_i_163_, last_key_i_164_, last_key_i_165_, last_key_i_166_, last_key_i_167_, last_key_i_168_, last_key_i_169_, last_key_i_170_, last_key_i_171_, last_key_i_172_, last_key_i_173_, last_key_i_174_, last_key_i_175_, last_key_i_176_, last_key_i_177_, last_key_i_178_, last_key_i_179_, last_key_i_180_, last_key_i_181_, last_key_i_182_, last_key_i_183_, last_key_i_184_, last_key_i_185_, last_key_i_186_, last_key_i_187_, last_key_i_188_, last_key_i_189_, last_key_i_190_, last_key_i_191_, new_key_o_0_, new_key_o_1_, new_key_o_2_, new_key_o_3_, new_key_o_4_, new_key_o_5_, new_key_o_6_, new_key_o_7_, new_key_o_8_, new_key_o_9_, new_key_o_10_, new_key_o_11_, new_key_o_12_, new_key_o_13_, new_key_o_14_, new_key_o_15_, new_key_o_16_, new_key_o_17_, new_key_o_18_, new_key_o_19_, new_key_o_20_, new_key_o_21_, new_key_o_22_, new_key_o_23_, new_key_o_24_, new_key_o_25_, new_key_o_26_, new_key_o_27_, new_key_o_28_, new_key_o_29_, new_key_o_30_, new_key_o_31_, new_key_o_32_, new_key_o_33_, new_key_o_34_, new_key_o_35_, new_key_o_36_, new_key_o_37_, new_key_o_38_, new_key_o_39_, new_key_o_40_, new_key_o_41_, new_key_o_42_, new_key_o_43_, new_key_o_44_, new_key_o_45_, new_key_o_46_, new_key_o_47_, new_key_o_48_, new_key_o_49_, new_key_o_50_, new_key_o_51_, new_key_o_52_, new_key_o_53_, new_key_o_54_, new_key_o_55_, new_key_o_56_, new_key_o_57_, new_key_o_58_, new_key_o_59_, new_key_o_60_, new_key_o_61_, new_key_o_62_, new_key_o_63_, new_key_o_64_, new_key_o_65_, new_key_o_66_, new_key_o_67_, new_key_o_68_, new_key_o_69_, new_key_o_70_, new_key_o_71_, new_key_o_72_, new_key_o_73_, new_key_o_74_, new_key_o_75_, new_key_o_76_, new_key_o_77_, new_key_o_78_, new_key_o_79_, new_key_o_80_, new_key_o_81_, new_key_o_82_, new_key_o_83_, new_key_o_84_, new_key_o_85_, new_key_o_86_, new_key_o_87_, new_key_o_88_, new_key_o_89_, new_key_o_90_, new_key_o_91_, new_key_o_92_, new_key_o_93_, new_key_o_94_, new_key_o_95_, new_key_o_96_, new_key_o_97_, new_key_o_98_, new_key_o_99_, new_key_o_100_, new_key_o_101_, new_key_o_102_, new_key_o_103_, new_key_o_104_, new_key_o_105_, new_key_o_106_, new_key_o_107_, new_key_o_108_, new_key_o_109_, new_key_o_110_, new_key_o_111_, new_key_o_112_, new_key_o_113_, new_key_o_114_, new_key_o_115_, new_key_o_116_, new_key_o_117_, new_key_o_118_, new_key_o_119_, new_key_o_120_, new_key_o_121_, new_key_o_122_, new_key_o_123_, new_key_o_124_, new_key_o_125_, new_key_o_126_, new_key_o_127_, new_key_o_128_, new_key_o_129_, new_key_o_130_, new_key_o_131_, new_key_o_132_, new_key_o_133_, new_key_o_134_, new_key_o_135_, new_key_o_136_, new_key_o_137_, new_key_o_138_, new_key_o_139_, new_key_o_140_, new_key_o_141_, new_key_o_142_, new_key_o_143_, new_key_o_144_, new_key_o_145_, new_key_o_146_, new_key_o_147_, new_key_o_148_, new_key_o_149_, new_key_o_150_, new_key_o_151_, new_key_o_152_, new_key_o_153_, new_key_o_154_, new_key_o_155_, new_key_o_156_, new_key_o_157_, new_key_o_158_, new_key_o_159_, new_key_o_160_, new_key_o_161_, new_key_o_162_, new_key_o_163_, new_key_o_164_, new_key_o_165_, new_key_o_166_, new_key_o_167_, new_key_o_168_, new_key_o_169_, new_key_o_170_, new_key_o_171_, new_key_o_172_, new_key_o_173_, new_key_o_174_, new_key_o_175_, new_key_o_176_, new_key_o_177_, new_key_o_178_, new_key_o_179_, new_key_o_180_, new_key_o_181_, new_key_o_182_, new_key_o_183_, new_key_o_184_, new_key_o_185_, new_key_o_186_, new_key_o_187_, new_key_o_188_, new_key_o_189_, new_key_o_190_, new_key_o_191_, ready_o, reset, round_i_0_, round_i_1_, round_i_2_, round_i_3_, sbox_access_o, sbox_data_i_0_, sbox_data_i_1_, sbox_data_i_2_, sbox_data_i_3_, sbox_data_i_4_, sbox_data_i_5_, sbox_data_i_6_, sbox_data_i_7_, sbox_data_o_0_, sbox_data_o_1_, sbox_data_o_2_, sbox_data_o_3_, sbox_data_o_4_, sbox_data_o_5_, sbox_data_o_6_, sbox_data_o_7_, sbox_decrypt_o, start_i);
input clk, last_key_i_0_, last_key_i_1_, last_key_i_2_, last_key_i_3_, last_key_i_4_, last_key_i_5_, last_key_i_6_, last_key_i_7_, last_key_i_8_, last_key_i_9_, last_key_i_10_, last_key_i_11_, last_key_i_12_, last_key_i_13_, last_key_i_14_, last_key_i_15_, last_key_i_16_, last_key_i_17_, last_key_i_18_, last_key_i_19_, last_key_i_20_, last_key_i_21_, last_key_i_22_, last_key_i_23_, last_key_i_24_, last_key_i_25_, last_key_i_26_, last_key_i_27_, last_key_i_28_, last_key_i_29_, last_key_i_30_, last_key_i_31_, last_key_i_32_, last_key_i_33_, last_key_i_34_, last_key_i_35_, last_key_i_36_, last_key_i_37_, last_key_i_38_, last_key_i_39_, last_key_i_40_, last_key_i_41_, last_key_i_42_, last_key_i_43_, last_key_i_44_, last_key_i_45_, last_key_i_46_, last_key_i_47_, last_key_i_48_, last_key_i_49_, last_key_i_50_, last_key_i_51_, last_key_i_52_, last_key_i_53_, last_key_i_54_, last_key_i_55_, last_key_i_56_, last_key_i_57_, last_key_i_58_, last_key_i_59_, last_key_i_60_, last_key_i_61_, last_key_i_62_, last_key_i_63_, last_key_i_64_, last_key_i_65_, last_key_i_66_, last_key_i_67_, last_key_i_68_, last_key_i_69_, last_key_i_70_, last_key_i_71_, last_key_i_72_, last_key_i_73_, last_key_i_74_, last_key_i_75_, last_key_i_76_, last_key_i_77_, last_key_i_78_, last_key_i_79_, last_key_i_80_, last_key_i_81_, last_key_i_82_, last_key_i_83_, last_key_i_84_, last_key_i_85_, last_key_i_86_, last_key_i_87_, last_key_i_88_, last_key_i_89_, last_key_i_90_, last_key_i_91_, last_key_i_92_, last_key_i_93_, last_key_i_94_, last_key_i_95_, last_key_i_96_, last_key_i_97_, last_key_i_98_, last_key_i_99_, last_key_i_100_, last_key_i_101_, last_key_i_102_, last_key_i_103_, last_key_i_104_, last_key_i_105_, last_key_i_106_, last_key_i_107_, last_key_i_108_, last_key_i_109_, last_key_i_110_, last_key_i_111_, last_key_i_112_, last_key_i_113_, last_key_i_114_, last_key_i_115_, last_key_i_116_, last_key_i_117_, last_key_i_118_, last_key_i_119_, last_key_i_120_, last_key_i_121_, last_key_i_122_, last_key_i_123_, last_key_i_124_, last_key_i_125_, last_key_i_126_, last_key_i_127_, last_key_i_128_, last_key_i_129_, last_key_i_130_, last_key_i_131_, last_key_i_132_, last_key_i_133_, last_key_i_134_, last_key_i_135_, last_key_i_136_, last_key_i_137_, last_key_i_138_, last_key_i_139_, last_key_i_140_, last_key_i_141_, last_key_i_142_, last_key_i_143_, last_key_i_144_, last_key_i_145_, last_key_i_146_, last_key_i_147_, last_key_i_148_, last_key_i_149_, last_key_i_150_, last_key_i_151_, last_key_i_152_, last_key_i_153_, last_key_i_154_, last_key_i_155_, last_key_i_156_, last_key_i_157_, last_key_i_158_, last_key_i_159_, last_key_i_160_, last_key_i_161_, last_key_i_162_, last_key_i_163_, last_key_i_164_, last_key_i_165_, last_key_i_166_, last_key_i_167_, last_key_i_168_, last_key_i_169_, last_key_i_170_, last_key_i_171_, last_key_i_172_, last_key_i_173_, last_key_i_174_, last_key_i_175_, last_key_i_176_, last_key_i_177_, last_key_i_178_, last_key_i_179_, last_key_i_180_, last_key_i_181_, last_key_i_182_, last_key_i_183_, last_key_i_184_, last_key_i_185_, last_key_i_186_, last_key_i_187_, last_key_i_188_, last_key_i_189_, last_key_i_190_, last_key_i_191_, reset, round_i_0_, round_i_1_, round_i_2_, round_i_3_, sbox_data_i_0_, sbox_data_i_1_, sbox_data_i_2_, sbox_data_i_3_, sbox_data_i_4_, sbox_data_i_5_, sbox_data_i_6_, sbox_data_i_7_, start_i;
output new_key_o_0_, new_key_o_1_, new_key_o_2_, new_key_o_3_, new_key_o_4_, new_key_o_5_, new_key_o_6_, new_key_o_7_, new_key_o_8_, new_key_o_9_, new_key_o_10_, new_key_o_11_, new_key_o_12_, new_key_o_13_, new_key_o_14_, new_key_o_15_, new_key_o_16_, new_key_o_17_, new_key_o_18_, new_key_o_19_, new_key_o_20_, new_key_o_21_, new_key_o_22_, new_key_o_23_, new_key_o_24_, new_key_o_25_, new_key_o_26_, new_key_o_27_, new_key_o_28_, new_key_o_29_, new_key_o_30_, new_key_o_31_, new_key_o_32_, new_key_o_33_, new_key_o_34_, new_key_o_35_, new_key_o_36_, new_key_o_37_, new_key_o_38_, new_key_o_39_, new_key_o_40_, new_key_o_41_, new_key_o_42_, new_key_o_43_, new_key_o_44_, new_key_o_45_, new_key_o_46_, new_key_o_47_, new_key_o_48_, new_key_o_49_, new_key_o_50_, new_key_o_51_, new_key_o_52_, new_key_o_53_, new_key_o_54_, new_key_o_55_, new_key_o_56_, new_key_o_57_, new_key_o_58_, new_key_o_59_, new_key_o_60_, new_key_o_61_, new_key_o_62_, new_key_o_63_, new_key_o_64_, new_key_o_65_, new_key_o_66_, new_key_o_67_, new_key_o_68_, new_key_o_69_, new_key_o_70_, new_key_o_71_, new_key_o_72_, new_key_o_73_, new_key_o_74_, new_key_o_75_, new_key_o_76_, new_key_o_77_, new_key_o_78_, new_key_o_79_, new_key_o_80_, new_key_o_81_, new_key_o_82_, new_key_o_83_, new_key_o_84_, new_key_o_85_, new_key_o_86_, new_key_o_87_, new_key_o_88_, new_key_o_89_, new_key_o_90_, new_key_o_91_, new_key_o_92_, new_key_o_93_, new_key_o_94_, new_key_o_95_, new_key_o_96_, new_key_o_97_, new_key_o_98_, new_key_o_99_, new_key_o_100_, new_key_o_101_, new_key_o_102_, new_key_o_103_, new_key_o_104_, new_key_o_105_, new_key_o_106_, new_key_o_107_, new_key_o_108_, new_key_o_109_, new_key_o_110_, new_key_o_111_, new_key_o_112_, new_key_o_113_, new_key_o_114_, new_key_o_115_, new_key_o_116_, new_key_o_117_, new_key_o_118_, new_key_o_119_, new_key_o_120_, new_key_o_121_, new_key_o_122_, new_key_o_123_, new_key_o_124_, new_key_o_125_, new_key_o_126_, new_key_o_127_, new_key_o_128_, new_key_o_129_, new_key_o_130_, new_key_o_131_, new_key_o_132_, new_key_o_133_, new_key_o_134_, new_key_o_135_, new_key_o_136_, new_key_o_137_, new_key_o_138_, new_key_o_139_, new_key_o_140_, new_key_o_141_, new_key_o_142_, new_key_o_143_, new_key_o_144_, new_key_o_145_, new_key_o_146_, new_key_o_147_, new_key_o_148_, new_key_o_149_, new_key_o_150_, new_key_o_151_, new_key_o_152_, new_key_o_153_, new_key_o_154_, new_key_o_155_, new_key_o_156_, new_key_o_157_, new_key_o_158_, new_key_o_159_, new_key_o_160_, new_key_o_161_, new_key_o_162_, new_key_o_163_, new_key_o_164_, new_key_o_165_, new_key_o_166_, new_key_o_167_, new_key_o_168_, new_key_o_169_, new_key_o_170_, new_key_o_171_, new_key_o_172_, new_key_o_173_, new_key_o_174_, new_key_o_175_, new_key_o_176_, new_key_o_177_, new_key_o_178_, new_key_o_179_, new_key_o_180_, new_key_o_181_, new_key_o_182_, new_key_o_183_, new_key_o_184_, new_key_o_185_, new_key_o_186_, new_key_o_187_, new_key_o_188_, new_key_o_189_, new_key_o_190_, new_key_o_191_, ready_o, sbox_access_o, sbox_data_o_0_, sbox_data_o_1_, sbox_data_o_2_, sbox_data_o_3_, sbox_data_o_4_, sbox_data_o_5_, sbox_data_o_6_, sbox_data_o_7_, sbox_decrypt_o;

sg13g2_nand3_1 U1 (.A(n36), .B(n826), .C(n37), .Y(sbox_data_o_1_));
sg13g2_nand3_1 U2 (.A(n26), .B(n985), .C(n27), .Y(sbox_data_o_3_));
sg13g2_o21ai_1 U3 (.A1(net25105), .A2(n226), .B1(n227), .Y(n767));
sg13g2_xnor2_1 U4 (.A(n153), .B(net25831), .Y(n154));
sg13g2_xnor2_1 U5 (.A(n537), .B(n803), .Y(n539));
sg13g2_inv_4 U6 (.A(last_key_i_1_), .Y(n39));
sg13g2_inv_4 U7 (.A(n854), .Y(n43));
sg13g2_inv_4 U8 (.A(last_key_i_11_), .Y(n864));
sg13g2_inv_4 U9 (.A(n827), .Y(n20));
sg13g2_inv_4 U10 (.A(n20), .Y(n25));
sg13g2_inv_4 U11 (.A(sbox_data_i_4_), .Y(n827));
sg13g2_inv_4 U12 (.A(n562), .Y(n563));
sg13g2_xnor2_1 U13 (.A(n565), .B(last_key_i_151_), .Y(n562));
sg13g2_o21ai_1 U14 (.A1(n807), .A2(net25107), .B1(n555), .Y(n699));
sg13g2_xnor2_1 U15 (.A(last_key_i_128_), .B(n347), .Y(n344));
sg13g2_o21ai_1 U16 (.A1(n337), .A2(net25097), .B1(n338), .Y(n609));
sg13g2_xnor2_1 U17 (.A(n44), .B(n335), .Y(n337));
sg13g2_o21ai_1 U18 (.A1(n539), .A2(net25109), .B1(n540), .Y(n693));
sg13g2_nand2_2 U19 (.A(last_key_i_91_), .B(n98), .Y(n975));
sg13g2_inv_4 U20 (.A(n98), .Y(n99));
sg13g2_buf_8 U21 (.A(last_key_i_133_), .X(n40));
sg13g2_xnor2_1 U22 (.A(last_key_i_123_), .B(n101), .Y(n98));
sg13g2_xnor2_1 U23 (.A(last_key_i_47_), .B(n190), .Y(n212));
sg13g2_nand2_2 U24 (.A(n282), .B(last_key_i_140_), .Y(n852));
sg13g2_xnor2_1 U25 (.A(last_key_i_164_), .B(col_4), .Y(n403));
sg13g2_nand2_2 U26 (.A(last_key_i_18_), .B(n9), .Y(n31));
sg13g2_xnor2_1 U27 (.A(last_key_i_132_), .B(n403), .Y(n400));
sg13g2_nand3_1 U28 (.A(n829), .B(n830), .C(n851), .Y(n853));
sg13g2_xnor2_1 U29 (.A(n54), .B(last_key_i_25_), .Y(n55));
sg13g2_xnor2_1 U30 (.A(last_key_i_57_), .B(n57), .Y(n54));
sg13g2_o21ai_1 U31 (.A1(n55), .A2(net25077), .B1(n56), .Y(n711));
sg13g2_inv_4 U32 (.A(n819), .Y(n46));
sg13g2_inv_4 U33 (.A(n46), .Y(n79));
sg13g2_o21ai_1 U34 (.A1(net25115), .A2(n276), .B1(n294), .Y(n794));
sg13g2_xnor2_1 U35 (.A(n115), .B(sbox_data_i_6_), .Y(n288));
sg13g2_xnor2_1 U36 (.A(n906), .B(n492), .Y(n496));
sg13g2_inv_4 U37 (.A(n800), .Y(n47));
sg13g2_inv_4 U38 (.A(n48), .Y(next_ready_o));
sg13g2_nand3_1 U39 (.A(n49), .B(n50), .C(state_2_), .Y(n48));
sg13g2_o21ai_1 U40 (.A1(n51), .A2(net25107), .B1(n53), .Y(n710));
sg13g2_nand2_2 U41 (.A(new_key_o_57_), .B(net25097), .Y(n53));
sg13g2_inv_4 U42 (.A(n54), .Y(n51));
sg13g2_o21ai_1 U43 (.A1(n494), .A2(net25111), .B1(n495), .Y(n675));
sg13g2_nand2_2 U44 (.A(new_key_o_25_), .B(net25083), .Y(n56));
sg13g2_inv_4 U45 (.A(n496), .Y(n494));
sg13g2_inv_4 U46 (.A(round_i_0_), .Y(n88));
sg13g2_o21ai_1 U47 (.A1(n57), .A2(net25105), .B1(n58), .Y(n712));
sg13g2_nand2_2 U48 (.A(new_key_o_89_), .B(net25107), .Y(n58));
sg13g2_nand2_2 U49 (.A(n88), .B(round_i_1_), .Y(n865));
sg13g2_o21ai_1 U50 (.A1(n60), .A2(net25105), .B1(n61), .Y(n713));
sg13g2_nand2_2 U51 (.A(new_key_o_121_), .B(net25097), .Y(n61));
sg13g2_inv_4 U52 (.A(n59), .Y(n60));
sg13g2_o21ai_1 U53 (.A1(net25103), .A2(n216), .B1(n217), .Y(n762));
sg13g2_o21ai_1 U54 (.A1(n62), .A2(net25105), .B1(n63), .Y(n714));
sg13g2_nand2_2 U55 (.A(new_key_o_153_), .B(net25093), .Y(n63));
sg13g2_xnor2_1 U56 (.A(n15), .B(n216), .Y(n234));
sg13g2_o21ai_1 U57 (.A1(n65), .A2(net25103), .B1(n66), .Y(n715));
sg13g2_nand2_2 U58 (.A(new_key_o_185_), .B(net25079), .Y(n66));
sg13g2_inv_4 U59 (.A(n64), .Y(n65));
sg13g2_inv_4 U60 (.A(n113), .Y(n115));
sg13g2_inv_4 U61 (.A(last_key_i_174_), .Y(n113));
sg13g2_o21ai_1 U62 (.A1(round_i_0_), .A2(n69), .B1(n70), .Y(n67));
sg13g2_o21ai_1 U63 (.A1(n243), .A2(net25105), .B1(n244), .Y(n773));
sg13g2_nand2_2 U64 (.A(new_key_o_58_), .B(net25075), .Y(n72));
sg13g2_nand2_2 U65 (.A(n312), .B(last_key_i_141_), .Y(n481));
sg13g2_nand2_2 U66 (.A(n892), .B(n891), .Y(n312));
sg13g2_nand2_2 U67 (.A(new_key_o_26_), .B(net25083), .Y(n75));
sg13g2_xnor2_1 U68 (.A(n409), .B(last_key_i_37_), .Y(n405));
sg13g2_inv_4 U69 (.A(n109), .Y(n186));
sg13g2_o21ai_1 U70 (.A1(n393), .A2(net25105), .B1(n394), .Y(n633));
sg13g2_nand2_2 U71 (.A(new_key_o_90_), .B(net25109), .Y(n77));
sg13g2_xnor2_1 U72 (.A(n24), .B(n391), .Y(n393));
sg13g2_o21ai_1 U73 (.A1(net25093), .A2(n945), .B1(n80), .Y(n719));
sg13g2_nand2_2 U74 (.A(new_key_o_122_), .B(net25081), .Y(n80));
sg13g2_o21ai_1 U75 (.A1(net25103), .A2(n220), .B1(n221), .Y(n764));
sg13g2_nand2_2 U76 (.A(n817), .B(last_key_i_136_), .Y(n845));
sg13g2_o21ai_1 U77 (.A1(net25115), .A2(n81), .B1(n82), .Y(n720));
sg13g2_nand2_2 U78 (.A(new_key_o_154_), .B(net25079), .Y(n82));
sg13g2_xnor2_1 U79 (.A(n83), .B(last_key_i_154_), .Y(n81));
sg13g2_o21ai_1 U80 (.A1(net25083), .A2(n84), .B1(n85), .Y(n721));
sg13g2_nand2_2 U81 (.A(new_key_o_186_), .B(net25111), .Y(n85));
sg13g2_inv_4 U82 (.A(n83), .Y(n84));
sg13g2_xnor2_1 U83 (.A(last_key_i_183_), .B(col_23_), .Y(n565));
sg13g2_xnor2_1 U84 (.A(last_key_i_159_), .B(n182), .Y(n179));
sg13g2_nor2_2 U85 (.A(n19), .B(n7), .Y(n18));
sg13g2_inv_4 U86 (.A(n856), .Y(n23));
sg13g2_inv_4 U87 (.A(last_key_i_172_), .Y(n828));
sg13g2_nand2_2 U88 (.A(new_key_o_59_), .B(net25113), .Y(n92));
sg13g2_xnor2_1 U89 (.A(n445), .B(last_key_i_135_), .Y(n442));
sg13g2_inv_4 U90 (.A(n804), .Y(n923));
sg13g2_nand2_2 U91 (.A(new_key_o_27_), .B(net25083), .Y(n95));
sg13g2_xnor2_1 U92 (.A(n431), .B(last_key_i_134_), .Y(n428));
sg13g2_inv_4 U93 (.A(last_key_i_173_), .Y(n890));
sg13g2_o21ai_1 U94 (.A1(net25109), .A2(n96), .B1(n97), .Y(n724));
sg13g2_nand2_2 U95 (.A(new_key_o_91_), .B(net25079), .Y(n97));
sg13g2_xnor2_1 U96 (.A(last_key_i_131_), .B(n389), .Y(n386));
sg13g2_o21ai_1 U97 (.A1(net25107), .A2(n99), .B1(n100), .Y(n725));
sg13g2_nand2_2 U98 (.A(new_key_o_123_), .B(net25093), .Y(n100));
sg13g2_xnor2_1 U99 (.A(n442), .B(last_key_i_103_), .Y(n440));
sg13g2_xnor2_1 U100 (.A(last_key_i_177_), .B(col_17_), .Y(n475));
sg13g2_o21ai_1 U101 (.A1(net25093), .A2(n101), .B1(n102), .Y(n726));
sg13g2_nand2_2 U102 (.A(new_key_o_155_), .B(net25093), .Y(n102));
sg13g2_xnor2_1 U103 (.A(last_key_i_179_), .B(col_19_), .Y(n505));
sg13g2_o21ai_1 U104 (.A1(net25103), .A2(n104), .B1(n105), .Y(n727));
sg13g2_nand2_2 U105 (.A(new_key_o_187_), .B(net25093), .Y(n105));
sg13g2_inv_4 U106 (.A(n103), .Y(n104));
sg13g2_inv_4 U107 (.A(n527), .Y(n929));
sg13g2_inv_4 U108 (.A(last_key_i_171_), .Y(n898));
sg13g2_inv_4 U109 (.A(last_key_i_140_), .Y(n851));
sg13g2_nand3_1 U110 (.A(n88), .B(n111), .C(n112), .Y(n108));
sg13g2_o21ai_1 U111 (.A1(net25105), .A2(n973), .B1(n114), .Y(n728));
sg13g2_nand2_2 U112 (.A(new_key_o_60_), .B(net25103), .Y(n114));
sg13g2_inv_4 U113 (.A(last_key_i_74_), .Y(n835));
sg13g2_o21ai_1 U114 (.A1(net25097), .A2(n116), .B1(n117), .Y(n729));
sg13g2_nand2_2 U115 (.A(new_key_o_28_), .B(net25077), .Y(n117));
sg13g2_xnor2_1 U116 (.A(n518), .B(n805), .Y(n116));
sg13g2_inv_4 U117 (.A(last_key_i_75_), .Y(n893));
sg13g2_o21ai_1 U118 (.A1(net25113), .A2(n118), .B1(n119), .Y(n730));
sg13g2_nand2_2 U119 (.A(new_key_o_92_), .B(net25097), .Y(n119));
sg13g2_o21ai_1 U120 (.A1(n228), .A2(net25105), .B1(n229), .Y(n768));
sg13g2_o21ai_1 U121 (.A1(net25077), .A2(n121), .B1(n122), .Y(n731));
sg13g2_nand2_2 U122 (.A(new_key_o_124_), .B(net25097), .Y(n122));
sg13g2_inv_4 U123 (.A(n120), .Y(n121));
sg13g2_nand2_2 U124 (.A(n866), .B(n131), .Y(n89));
sg13g2_o21ai_1 U125 (.A1(net25093), .A2(n123), .B1(n124), .Y(n732));
sg13g2_nand2_2 U126 (.A(new_key_o_156_), .B(net25097), .Y(n124));
sg13g2_inv_4 U127 (.A(n865), .Y(n866));
sg13g2_o21ai_1 U128 (.A1(net25111), .A2(n126), .B1(n127), .Y(n733));
sg13g2_nand2_2 U129 (.A(new_key_o_188_), .B(net25093), .Y(n127));
sg13g2_inv_4 U130 (.A(n125), .Y(n126));
sg13g2_nand2_2 U131 (.A(n914), .B(n913), .Y(n916));
sg13g2_inv_4 U132 (.A(n487), .Y(n914));
sg13g2_nand2_2 U133 (.A(n932), .B(n931), .Y(n934));
sg13g2_nand2_2 U134 (.A(n949), .B(n948), .Y(n951));
sg13g2_nand2_2 U135 (.A(n112), .B(n132), .Y(n130));
sg13g2_o21ai_1 U136 (.A1(net25113), .A2(n962), .B1(n134), .Y(n734));
sg13g2_nand2_2 U137 (.A(new_key_o_61_), .B(net25079), .Y(n134));
sg13g2_nand2_2 U138 (.A(n438), .B(n868), .Y(n870));
sg13g2_o21ai_1 U139 (.A1(last_key_i_87_), .A2(n560), .B1(n860), .Y(n557));
sg13g2_nand2_2 U140 (.A(new_key_o_29_), .B(net25093), .Y(n137));
sg13g2_nand3_1 U141 (.A(n50), .B(n318), .C(state_0_), .Y(n45));
sg13g2_nand2_2 U142 (.A(n918), .B(n917), .Y(n920));
sg13g2_o21ai_1 U143 (.A1(net25111), .A2(n138), .B1(n139), .Y(n736));
sg13g2_nand2_2 U144 (.A(new_key_o_93_), .B(net25127), .Y(n139));
sg13g2_nand2_2 U145 (.A(n940), .B(n939), .Y(n942));
sg13g2_o21ai_1 U146 (.A1(net25113), .A2(n141), .B1(n142), .Y(n737));
sg13g2_nand2_2 U147 (.A(new_key_o_125_), .B(net25103), .Y(n142));
sg13g2_inv_4 U148 (.A(n140), .Y(n141));
sg13g2_inv_4 U149 (.A(n520), .Y(n940));
sg13g2_o21ai_1 U150 (.A1(net25097), .A2(n143), .B1(n144), .Y(n738));
sg13g2_nand2_2 U151 (.A(new_key_o_157_), .B(net25097), .Y(n144));
sg13g2_nand2_2 U152 (.A(n373), .B(n526), .Y(n541));
sg13g2_o21ai_1 U153 (.A1(net25115), .A2(n146), .B1(n147), .Y(n739));
sg13g2_nand2_2 U154 (.A(new_key_o_189_), .B(net25093), .Y(n147));
sg13g2_inv_4 U155 (.A(n145), .Y(n146));
sg13g2_o21ai_1 U156 (.A1(last_key_i_53_), .A2(n527), .B1(n930), .Y(n522));
sg13g2_o21ai_1 U157 (.A1(last_key_i_86_), .A2(n545), .B1(n900), .Y(n542));
sg13g2_nand2_2 U158 (.A(n945), .B(n944), .Y(n947));
sg13g2_nand3_1 U159 (.A(round_i_1_), .B(n88), .C(n112), .Y(n150));
sg13g2_inv_4 U160 (.A(n78), .Y(n945));
sg13g2_nand2_2 U161 (.A(n959), .B(n958), .Y(n961));
sg13g2_nand2_2 U162 (.A(new_key_o_62_), .B(net25127), .Y(n152));
sg13g2_inv_4 U163 (.A(n153), .Y(n151));
sg13g2_nand2_2 U164 (.A(n285), .B(n270), .Y(n306));
sg13g2_nand2_2 U165 (.A(new_key_o_30_), .B(net25083), .Y(n155));
sg13g2_nand2_2 U166 (.A(n836), .B(n835), .Y(n838));
sg13g2_nand3_1 U167 (.A(n49), .B(n318), .C(state_1_), .Y(n1));
sg13g2_o21ai_1 U168 (.A1(net25115), .A2(n156), .B1(n157), .Y(n742));
sg13g2_nand2_2 U169 (.A(new_key_o_94_), .B(net25107), .Y(n157));
sg13g2_nand3_1 U170 (.A(n21), .B(n986), .C(n22), .Y(sbox_data_o_4_));
sg13g2_o21ai_1 U171 (.A1(net25115), .A2(n159), .B1(n160), .Y(n743));
sg13g2_nand2_2 U172 (.A(new_key_o_126_), .B(net25081), .Y(n160));
sg13g2_inv_4 U173 (.A(n158), .Y(n159));
sg13g2_nand3_1 U174 (.A(n42), .B(n987), .C(n41), .Y(sbox_data_o_0_));
sg13g2_o21ai_1 U175 (.A1(net25115), .A2(n161), .B1(n162), .Y(n744));
sg13g2_nand2_2 U176 (.A(new_key_o_158_), .B(net25097), .Y(n162));
sg13g2_nand2_2 U177 (.A(n524), .B(n433), .Y(n867));
sg13g2_o21ai_1 U178 (.A1(net25079), .A2(n164), .B1(n165), .Y(n745));
sg13g2_nand2_2 U179 (.A(new_key_o_190_), .B(net25079), .Y(n165));
sg13g2_inv_4 U180 (.A(n163), .Y(n164));
sg13g2_o21ai_1 U181 (.A1(last_key_i_34_), .A2(n367), .B1(n887), .Y(n363));
sg13g2_o21ai_1 U182 (.A1(last_key_i_67_), .A2(n384), .B1(n878), .Y(n381));
sg13g2_nand2_2 U183 (.A(n429), .B(n871), .Y(n873));
sg13g2_nand3_1 U184 (.A(round_i_0_), .B(round_i_1_), .C(n112), .Y(n168));
sg13g2_o21ai_1 U185 (.A1(last_key_i_112_), .A2(n457), .B1(n921), .Y(n455));
sg13g2_o21ai_1 U186 (.A1(last_key_i_115_), .A2(n502), .B1(n908), .Y(n500));
sg13g2_nand2_2 U187 (.A(n936), .B(n935), .Y(n938));
sg13g2_nand2_2 U188 (.A(new_key_o_63_), .B(net25109), .Y(n170));
sg13g2_nand2_2 U189 (.A(n969), .B(n968), .Y(n971));
sg13g2_nand2_2 U190 (.A(new_key_o_31_), .B(net25093), .Y(n172));
sg13g2_inv_4 U191 (.A(n173), .Y(n171));
sg13g2_xnor2_1 U192 (.A(n106), .B(n107), .Y(n103));
sg13g2_o21ai_1 U193 (.A1(last_key_i_124_), .A2(n123), .B1(n972), .Y(n120));
sg13g2_o21ai_1 U194 (.A1(net25081), .A2(n175), .B1(n176), .Y(n748));
sg13g2_nand2_2 U195 (.A(new_key_o_95_), .B(net25075), .Y(n176));
sg13g2_nand3_1 U196 (.A(n460), .B(n891), .C(n892), .Y(n488));
sg13g2_o21ai_1 U197 (.A1(n952), .A2(n45), .B1(n305), .Y(n585));
sg13g2_o21ai_1 U198 (.A1(net25075), .A2(n177), .B1(n178), .Y(n749));
sg13g2_nand2_2 U199 (.A(new_key_o_127_), .B(net25097), .Y(n178));
sg13g2_o21ai_1 U200 (.A1(n524), .A2(n433), .B1(n867), .Y(n435));
sg13g2_o21ai_1 U201 (.A1(net25075), .A2(n180), .B1(n181), .Y(n750));
sg13g2_nand2_2 U202 (.A(new_key_o_159_), .B(net25103), .Y(n181));
sg13g2_inv_4 U203 (.A(n179), .Y(n180));
sg13g2_xnor2_1 U204 (.A(n977), .B(n477), .Y(n479));
sg13g2_o21ai_1 U205 (.A1(net25127), .A2(n182), .B1(n183), .Y(n751));
sg13g2_nand2_2 U206 (.A(new_key_o_191_), .B(net25083), .Y(n183));
sg13g2_xnor2_1 U207 (.A(n926), .B(n522), .Y(n806));
sg13g2_xnor2_1 U208 (.A(n552), .B(net25888), .Y(n807));
sg13g2_nand3_1 U209 (.A(n3), .B(n988), .C(n4), .Y(sbox_data_o_7_));
sg13g2_xnor2_1 U210 (.A(n978), .B(n567), .Y(n569));
sg13g2_xnor2_1 U211 (.A(n979), .B(n962), .Y(n136));
sg13g2_xnor2_1 U212 (.A(n30), .B(n222), .Y(n243));
sg13g2_xnor2_1 U213 (.A(n2), .B(n212), .Y(n228));
sg13g2_nand2_2 U214 (.A(n230), .B(last_key_i_79_), .Y(n253));
sg13g2_o21ai_1 U215 (.A1(n188), .A2(net25103), .B1(n189), .Y(n752));
sg13g2_nand2_2 U216 (.A(new_key_o_79_), .B(net25127), .Y(n189));
sg13g2_inv_4 U217 (.A(n190), .Y(n188));
sg13g2_o21ai_1 U218 (.A1(n191), .A2(net25127), .B1(n192), .Y(n753));
sg13g2_nand2_2 U219 (.A(new_key_o_78_), .B(net25103), .Y(n192));
sg13g2_inv_4 U220 (.A(n193), .Y(n191));
sg13g2_o21ai_1 U221 (.A1(n194), .A2(net25127), .B1(n195), .Y(n754));
sg13g2_nand2_2 U222 (.A(new_key_o_77_), .B(net25075), .Y(n195));
sg13g2_nand2_2 U223 (.A(n133), .B(n135), .Y(n261));
sg13g2_o21ai_1 U224 (.A1(n197), .A2(net25103), .B1(n198), .Y(n755));
sg13g2_nand2_2 U225 (.A(new_key_o_76_), .B(net25075), .Y(n198));
sg13g2_inv_4 U226 (.A(n199), .Y(n197));
sg13g2_o21ai_1 U227 (.A1(n200), .A2(net25103), .B1(n201), .Y(n756));
sg13g2_nand2_2 U228 (.A(new_key_o_75_), .B(net25075), .Y(n201));
sg13g2_inv_4 U229 (.A(n202), .Y(n200));
sg13g2_o21ai_1 U230 (.A1(n203), .A2(net25103), .B1(n204), .Y(n757));
sg13g2_nand2_2 U231 (.A(new_key_o_74_), .B(net25075), .Y(n204));
sg13g2_inv_4 U232 (.A(n205), .Y(n203));
sg13g2_o21ai_1 U233 (.A1(net25103), .A2(n206), .B1(n207), .Y(n758));
sg13g2_nand2_2 U234 (.A(new_key_o_73_), .B(net25075), .Y(n207));
sg13g2_nand2_2 U235 (.A(n253), .B(n261), .Y(n190));
sg13g2_o21ai_1 U236 (.A1(n209), .A2(net25103), .B1(n210), .Y(n759));
sg13g2_nand2_2 U237 (.A(new_key_o_72_), .B(net25077), .Y(n210));
sg13g2_inv_4 U238 (.A(n211), .Y(n209));
sg13g2_inv_4 U239 (.A(n230), .Y(n133));
sg13g2_nand2_2 U240 (.A(new_key_o_47_), .B(net25077), .Y(n213));
sg13g2_inv_4 U241 (.A(last_key_i_79_), .Y(n135));
sg13g2_nand2_2 U242 (.A(new_key_o_46_), .B(net25077), .Y(n215));
sg13g2_nand2_2 U243 (.A(n291), .B(last_key_i_143_), .Y(n304));
sg13g2_nand2_2 U244 (.A(new_key_o_45_), .B(net25077), .Y(n217));
sg13g2_o21ai_1 U245 (.A1(net25105), .A2(n218), .B1(n219), .Y(n763));
sg13g2_nand2_2 U246 (.A(new_key_o_44_), .B(net25079), .Y(n219));
sg13g2_nand2_2 U247 (.A(n304), .B(n306), .Y(n267));
sg13g2_nand2_2 U248 (.A(new_key_o_43_), .B(net25079), .Y(n221));
sg13g2_inv_4 U249 (.A(last_key_i_143_), .Y(n270));
sg13g2_nand2_2 U250 (.A(new_key_o_42_), .B(net25079), .Y(n223));
sg13g2_inv_4 U251 (.A(n291), .Y(n285));
sg13g2_nand2_2 U252 (.A(new_key_o_41_), .B(net25081), .Y(n225));
sg13g2_inv_4 U253 (.A(n981), .Y(n308));
sg13g2_nand2_2 U254 (.A(new_key_o_40_), .B(net25081), .Y(n227));
sg13g2_xnor2_1 U255 (.A(last_key_i_175_), .B(sbox_data_i_7_), .Y(n291));
sg13g2_nand2_2 U256 (.A(new_key_o_15_), .B(net25081), .Y(n229));
sg13g2_inv_4 U257 (.A(n414), .Y(n310));
sg13g2_a21oi_2 U258 (.A1(net39266), .A2(last_key_i_24_), .B1(n43), .Y(n42));
sg13g2_nand2_2 U259 (.A(last_key_i_19_), .B(n9), .Y(n26));
sg13g2_xnor2_1 U260 (.A(last_key_i_168_), .B(sbox_data_i_0_), .Y(n817));
sg13g2_nand2_2 U261 (.A(n897), .B(n898), .Y(n808));
sg13g2_nand2_2 U262 (.A(new_key_o_14_), .B(net25081), .Y(n232));
sg13g2_xnor2_1 U263 (.A(n40), .B(n417), .Y(n904));
sg13g2_inv_4 U264 (.A(n372), .Y(n373));
sg13g2_xnor2_1 U265 (.A(last_key_i_176_), .B(col_16_), .Y(n804));
sg13g2_inv_4 U266 (.A(sbox_data_i_1_), .Y(n414));
sg13g2_inv_4 U267 (.A(n310), .Y(n952));
sg13g2_nand2_2 U268 (.A(new_key_o_13_), .B(net25083), .Y(n235));
sg13g2_nand2_2 U269 (.A(n481), .B(n488), .Y(n424));
sg13g2_xnor2_1 U270 (.A(last_key_i_166_), .B(col_6), .Y(n431));
sg13g2_xnor2_1 U271 (.A(n864), .B(n220), .Y(n240));
sg13g2_nand2_2 U272 (.A(n481), .B(n488), .Y(n263));
sg13g2_inv_4 U273 (.A(last_key_i_141_), .Y(n460));
sg13g2_nand2_2 U274 (.A(new_key_o_12_), .B(net25083), .Y(n238));
sg13g2_nand2_2 U275 (.A(last_key_i_21_), .B(n9), .Y(n16));
sg13g2_nand2_2 U276 (.A(last_key_i_20_), .B(n9), .Y(n21));
sg13g2_nand2_2 U277 (.A(n218), .B(n943), .Y(n888));
sg13g2_xnor2_1 U278 (.A(n467), .B(last_key_i_49_), .Y(n462));
sg13g2_xnor2_1 U279 (.A(last_key_i_81_), .B(n470), .Y(n467));
sg13g2_nand2_2 U280 (.A(new_key_o_11_), .B(net25083), .Y(n241));
sg13g2_inv_4 U281 (.A(last_key_i_12_), .Y(n943));
sg13g2_inv_4 U282 (.A(last_key_i_28_), .Y(n503));
sg13g2_inv_4 U283 (.A(n503), .Y(n518));
sg13g2_o21ai_1 U284 (.A1(net25105), .A2(n224), .B1(n225), .Y(n766));
sg13g2_xnor2_1 U285 (.A(last_key_i_167_), .B(col_7), .Y(n445));
sg13g2_nand2_2 U286 (.A(new_key_o_10_), .B(net25093), .Y(n244));
sg13g2_a21oi_2 U287 (.A1(last_key_i_25_), .A2(n5), .B1(n38), .Y(n37));
sg13g2_inv_4 U288 (.A(net39263), .Y(net39266));
sg13g2_nand3_1 U289 (.A(n16), .B(n989), .C(n17), .Y(sbox_data_o_5_));
sg13g2_nand4_1 U290 (.A(last_key_i_0_), .B(state_0_), .C(state_1_), .D(n318), .Y(n854));
sg13g2_inv_4 U291 (.A(net26231), .Y(n524));
sg13g2_nand2_2 U292 (.A(new_key_o_9_), .B(net25083), .Y(n247));
sg13g2_xnor2_1 U293 (.A(last_key_i_120_), .B(n577), .Y(n575));
sg13g2_nand2_2 U294 (.A(n372), .B(last_key_i_98_), .Y(n528));
sg13g2_nand2_2 U295 (.A(n528), .B(n541), .Y(n370));
sg13g2_inv_4 U296 (.A(last_key_i_98_), .Y(n526));
sg13g2_nand2_2 U297 (.A(n375), .B(last_key_i_130_), .Y(n571));
sg13g2_nand2_2 U298 (.A(new_key_o_8_), .B(net25083), .Y(n250));
sg13g2_nand2_2 U299 (.A(n554), .B(n556), .Y(n802));
sg13g2_nand2_2 U300 (.A(n571), .B(n802), .Y(n372));
sg13g2_inv_4 U301 (.A(n375), .Y(n554));
sg13g2_inv_4 U302 (.A(last_key_i_130_), .Y(n556));
sg13g2_o21ai_1 U303 (.A1(net25127), .A2(n251), .B1(n252), .Y(n776));
sg13g2_nand2_2 U304 (.A(new_key_o_104_), .B(net25083), .Y(n252));
sg13g2_xnor2_1 U305 (.A(n370), .B(last_key_i_66_), .Y(n367));
sg13g2_o21ai_1 U306 (.A1(net25127), .A2(n308), .B1(n254), .Y(n777));
sg13g2_nand2_2 U307 (.A(new_key_o_105_), .B(net25083), .Y(n254));
sg13g2_o21ai_1 U308 (.A1(net25111), .A2(n370), .B1(n371), .Y(n623));
sg13g2_o21ai_1 U309 (.A1(net25127), .A2(n245), .B1(n256), .Y(n778));
sg13g2_nand2_2 U310 (.A(new_key_o_106_), .B(net25083), .Y(n256));
sg13g2_inv_4 U311 (.A(last_key_i_22_), .Y(n803));
sg13g2_o21ai_1 U312 (.A1(net25127), .A2(n242), .B1(n258), .Y(n779));
sg13g2_nand2_2 U313 (.A(new_key_o_107_), .B(net25083), .Y(n258));
sg13g2_xnor2_1 U314 (.A(last_key_i_117_), .B(n532), .Y(n530));
sg13g2_o21ai_1 U315 (.A1(net25127), .A2(n239), .B1(n260), .Y(n780));
sg13g2_nand2_2 U316 (.A(new_key_o_108_), .B(net25083), .Y(n260));
sg13g2_xnor2_1 U317 (.A(last_key_i_149_), .B(n535), .Y(n532));
sg13g2_o21ai_1 U318 (.A1(net25127), .A2(n236), .B1(n262), .Y(n781));
sg13g2_nand2_2 U319 (.A(new_key_o_109_), .B(net25081), .Y(n262));
sg13g2_xnor2_1 U320 (.A(last_key_i_181_), .B(col_21_), .Y(n535));
sg13g2_o21ai_1 U321 (.A1(net25127), .A2(n233), .B1(n264), .Y(n782));
sg13g2_nand2_2 U322 (.A(new_key_o_110_), .B(net25081), .Y(n264));
sg13g2_inv_4 U323 (.A(last_key_i_8_), .Y(n984));
sg13g2_o21ai_1 U324 (.A1(n230), .A2(net25103), .B1(n266), .Y(n783));
sg13g2_nand2_2 U325 (.A(new_key_o_111_), .B(net25081), .Y(n266));
sg13g2_inv_4 U326 (.A(n502), .Y(n907));
sg13g2_o21ai_1 U327 (.A1(n268), .A2(net25115), .B1(n269), .Y(n784));
sg13g2_nand2_2 U328 (.A(new_key_o_136_), .B(net25081), .Y(n269));
sg13g2_inv_4 U329 (.A(n810), .Y(n268));
sg13g2_inv_4 U330 (.A(n517), .Y(n936));
sg13g2_o21ai_1 U331 (.A1(n271), .A2(net25083), .B1(n272), .Y(n785));
sg13g2_nand2_2 U332 (.A(new_key_o_137_), .B(net25081), .Y(n272));
sg13g2_inv_4 U333 (.A(n255), .Y(n271));
sg13g2_inv_4 U334 (.A(n5), .Y(net39263));
sg13g2_o21ai_1 U335 (.A1(n274), .A2(net25083), .B1(n275), .Y(n786));
sg13g2_nand2_2 U336 (.A(new_key_o_138_), .B(net25081), .Y(n275));
sg13g2_inv_4 U337 (.A(n257), .Y(n274));
sg13g2_nand2_2 U338 (.A(last_key_i_124_), .B(n123), .Y(n972));
sg13g2_o21ai_1 U339 (.A1(n277), .A2(net25079), .B1(n278), .Y(n787));
sg13g2_nand2_2 U340 (.A(new_key_o_139_), .B(net25081), .Y(n278));
sg13g2_inv_4 U341 (.A(n259), .Y(n277));
sg13g2_xnor2_1 U342 (.A(last_key_i_189_), .B(col_29_), .Y(n149));
sg13g2_o21ai_1 U343 (.A1(n280), .A2(net25109), .B1(n281), .Y(n788));
sg13g2_nand2_2 U344 (.A(new_key_o_140_), .B(net25079), .Y(n281));
sg13g2_inv_4 U345 (.A(n809), .Y(n280));
sg13g2_o21ai_1 U346 (.A1(n449), .A2(net25115), .B1(n450), .Y(n657));
sg13g2_o21ai_1 U347 (.A1(n283), .A2(net25097), .B1(n284), .Y(n789));
sg13g2_nand2_2 U348 (.A(new_key_o_141_), .B(net25079), .Y(n284));
sg13g2_inv_4 U349 (.A(n424), .Y(n283));
sg13g2_xnor2_1 U350 (.A(last_key_i_186_), .B(col_26_), .Y(n87));
sg13g2_o21ai_1 U351 (.A1(n286), .A2(net25093), .B1(n287), .Y(n790));
sg13g2_nand2_2 U352 (.A(new_key_o_142_), .B(net25079), .Y(n287));
sg13g2_inv_4 U353 (.A(n265), .Y(n286));
sg13g2_xnor2_1 U354 (.A(n86), .B(n87), .Y(n83));
sg13g2_o21ai_1 U355 (.A1(n289), .A2(net25127), .B1(n290), .Y(n791));
sg13g2_nand2_2 U356 (.A(new_key_o_143_), .B(net25079), .Y(n290));
sg13g2_inv_4 U357 (.A(n267), .Y(n289));
sg13g2_xnor2_1 U358 (.A(last_key_i_158_), .B(n163), .Y(n161));
sg13g2_o21ai_1 U359 (.A1(n817), .A2(net25077), .B1(n292), .Y(n792));
sg13g2_nand2_2 U360 (.A(new_key_o_168_), .B(net25079), .Y(n292));
sg13g2_xnor2_1 U361 (.A(last_key_i_92_), .B(n120), .Y(n118));
sg13g2_o21ai_1 U362 (.A1(net25107), .A2(n273), .B1(n293), .Y(n793));
sg13g2_nand2_2 U363 (.A(new_key_o_169_), .B(net25079), .Y(n293));
sg13g2_inv_4 U364 (.A(n805), .Y(n973));
sg13g2_o21ai_1 U365 (.A1(net25107), .A2(n151), .B1(n152), .Y(n740));
sg13g2_nand2_2 U366 (.A(new_key_o_170_), .B(net25079), .Y(n294));
sg13g2_nand2_2 U367 (.A(n852), .B(n853), .Y(n809));
sg13g2_xnor2_1 U368 (.A(n452), .B(last_key_i_48_), .Y(n447));
sg13g2_nand2_2 U369 (.A(new_key_o_171_), .B(net25079), .Y(n295));
sg13g2_xnor2_1 U370 (.A(last_key_i_60_), .B(n118), .Y(n805));
sg13g2_o21ai_1 U371 (.A1(n282), .A2(net25113), .B1(n296), .Y(n796));
sg13g2_nand2_2 U372 (.A(new_key_o_172_), .B(net25077), .Y(n296));
sg13g2_xnor2_1 U373 (.A(n128), .B(n129), .Y(n125));
sg13g2_xnor2_1 U374 (.A(last_key_i_157_), .B(n145), .Y(n143));
sg13g2_nand2_2 U375 (.A(new_key_o_173_), .B(net25077), .Y(n297));
sg13g2_xnor2_1 U376 (.A(last_key_i_187_), .B(col_27_), .Y(n107));
sg13g2_o21ai_1 U377 (.A1(net25079), .A2(n288), .B1(n298), .Y(n798));
sg13g2_nand2_2 U378 (.A(new_key_o_174_), .B(net25077), .Y(n298));
sg13g2_o21ai_1 U379 (.A1(net25079), .A2(n91), .B1(n92), .Y(n722));
sg13g2_o21ai_1 U380 (.A1(net25093), .A2(n291), .B1(n299), .Y(n799));
sg13g2_nand2_2 U381 (.A(new_key_o_175_), .B(net25077), .Y(n299));
sg13g2_inv_4 U382 (.A(n93), .Y(n91));
sg13g2_nand2_2 U383 (.A(n1), .B(n45), .Y(n800));
sg13g2_nand2_2 U384 (.A(net39263), .B(n1), .Y(n801));
sg13g2_xnor2_1 U385 (.A(n395), .B(last_key_i_36_), .Y(n391));
sg13g2_xnor2_1 U386 (.A(last_key_i_185_), .B(col_25_), .Y(n68));
sg13g2_inv_4 U387 (.A(start_i), .Y(n300));
sg13g2_o21ai_1 U388 (.A1(n45), .A2(n302), .B1(n303), .Y(n584));
sg13g2_nand2_2 U389 (.A(col_0), .B(n45), .Y(n303));
sg13g2_o21ai_1 U390 (.A1(n154), .A2(net25105), .B1(n155), .Y(n741));
sg13g2_nand2_2 U391 (.A(col_1), .B(n45), .Y(n305));
sg13g2_o21ai_1 U392 (.A1(n45), .A2(n79), .B1(n307), .Y(n586));
sg13g2_nand2_2 U393 (.A(col_2), .B(n45), .Y(n307));
sg13g2_o21ai_1 U394 (.A1(n45), .A2(n897), .B1(n309), .Y(n587));
sg13g2_nand2_2 U395 (.A(col_3), .B(n45), .Y(n309));
sg13g2_o21ai_1 U396 (.A1(n45), .A2(n25), .B1(n311), .Y(n588));
sg13g2_nand2_2 U397 (.A(col_4), .B(n45), .Y(n311));
sg13g2_o21ai_1 U398 (.A1(n45), .A2(n889), .B1(n313), .Y(n589));
sg13g2_nand2_2 U399 (.A(col_5), .B(n45), .Y(n313));
sg13g2_o21ai_1 U400 (.A1(n45), .A2(n314), .B1(n315), .Y(n590));
sg13g2_nand2_2 U401 (.A(col_6), .B(n45), .Y(n315));
sg13g2_o21ai_1 U402 (.A1(n45), .A2(n316), .B1(n317), .Y(n591));
sg13g2_nand2_2 U403 (.A(col_7), .B(n45), .Y(n317));
sg13g2_nand2_2 U404 (.A(n845), .B(n846), .Y(n810));
sg13g2_o21ai_1 U405 (.A1(n7), .A2(n302), .B1(n319), .Y(n592));
sg13g2_nand2_2 U406 (.A(col_16_), .B(n7), .Y(n319));
sg13g2_o21ai_1 U407 (.A1(n7), .A2(n952), .B1(n320), .Y(n593));
sg13g2_nand2_2 U408 (.A(col_17_), .B(n7), .Y(n320));
sg13g2_o21ai_1 U409 (.A1(n7), .A2(n79), .B1(n321), .Y(n594));
sg13g2_nand2_2 U410 (.A(col_18_), .B(n7), .Y(n321));
sg13g2_o21ai_1 U411 (.A1(n7), .A2(n897), .B1(n322), .Y(n595));
sg13g2_nand2_2 U412 (.A(col_19_), .B(n7), .Y(n322));
sg13g2_o21ai_1 U413 (.A1(n7), .A2(n25), .B1(n323), .Y(n596));
sg13g2_nand2_2 U414 (.A(col_20_), .B(n7), .Y(n323));
sg13g2_o21ai_1 U415 (.A1(n7), .A2(n889), .B1(n324), .Y(n597));
sg13g2_nand2_2 U416 (.A(col_21_), .B(n7), .Y(n324));
sg13g2_o21ai_1 U417 (.A1(n7), .A2(n314), .B1(n325), .Y(n598));
sg13g2_nand2_2 U418 (.A(col_22_), .B(n7), .Y(n325));
sg13g2_o21ai_1 U419 (.A1(n7), .A2(n316), .B1(n326), .Y(n599));
sg13g2_nand2_2 U420 (.A(col_23_), .B(n7), .Y(n326));
sg13g2_o21ai_1 U421 (.A1(n1), .A2(n302), .B1(n327), .Y(n600));
sg13g2_nand2_2 U422 (.A(col_24_), .B(n1), .Y(n327));
sg13g2_inv_4 U423 (.A(sbox_data_i_0_), .Y(n302));
sg13g2_o21ai_1 U424 (.A1(n1), .A2(n952), .B1(n328), .Y(n601));
sg13g2_nand2_2 U425 (.A(col_25_), .B(n1), .Y(n328));
sg13g2_xnor2_1 U426 (.A(n859), .B(n73), .Y(n74));
sg13g2_o21ai_1 U427 (.A1(n1), .A2(n79), .B1(n329), .Y(n602));
sg13g2_nand2_2 U428 (.A(col_26_), .B(n1), .Y(n329));
sg13g2_inv_4 U429 (.A(sbox_data_i_3_), .Y(n897));
sg13g2_o21ai_1 U430 (.A1(n1), .A2(n897), .B1(n330), .Y(n603));
sg13g2_nand2_2 U431 (.A(col_27_), .B(n1), .Y(n330));
sg13g2_o21ai_1 U432 (.A1(net25075), .A2(n71), .B1(n72), .Y(n716));
sg13g2_o21ai_1 U433 (.A1(n1), .A2(n25), .B1(n331), .Y(n604));
sg13g2_nand2_2 U434 (.A(col_28_), .B(n1), .Y(n331));
sg13g2_inv_4 U435 (.A(n73), .Y(n71));
sg13g2_o21ai_1 U436 (.A1(n1), .A2(n889), .B1(n332), .Y(n605));
sg13g2_nand2_2 U437 (.A(col_29_), .B(n1), .Y(n332));
sg13g2_o21ai_1 U438 (.A1(n569), .A2(net25107), .B1(n570), .Y(n705));
sg13g2_o21ai_1 U439 (.A1(n1), .A2(n314), .B1(n333), .Y(n606));
sg13g2_nand2_2 U440 (.A(col_30_), .B(n1), .Y(n333));
sg13g2_inv_4 U441 (.A(sbox_data_i_6_), .Y(n314));
sg13g2_o21ai_1 U442 (.A1(n1), .A2(n316), .B1(n334), .Y(n607));
sg13g2_nand2_2 U443 (.A(col_31_), .B(n1), .Y(n334));
sg13g2_inv_4 U444 (.A(sbox_data_i_7_), .Y(n316));
sg13g2_o21ai_1 U445 (.A1(n212), .A2(net25103), .B1(n213), .Y(n760));
sg13g2_o21ai_1 U446 (.A1(net25103), .A2(n335), .B1(n336), .Y(n608));
sg13g2_nand2_2 U447 (.A(new_key_o_32_), .B(net25077), .Y(n336));
sg13g2_xnor2_1 U448 (.A(last_key_i_190_), .B(col_30_), .Y(n167));
sg13g2_nand2_2 U449 (.A(new_key_o_0_), .B(net25077), .Y(n338));
sg13g2_a21oi_2 U450 (.A1(last_key_i_30_), .A2(n5), .B1(n13), .Y(n12));
sg13g2_o21ai_1 U451 (.A1(n222), .A2(net25103), .B1(n223), .Y(n765));
sg13g2_inv_4 U452 (.A(n208), .Y(n206));
sg13g2_o21ai_1 U453 (.A1(n340), .A2(net25075), .B1(n341), .Y(n610));
sg13g2_nand2_2 U454 (.A(new_key_o_64_), .B(net25077), .Y(n341));
sg13g2_inv_4 U455 (.A(n339), .Y(n340));
sg13g2_nand3_1 U456 (.A(n131), .B(round_i_1_), .C(round_i_0_), .Y(n110));
sg13g2_o21ai_1 U457 (.A1(n342), .A2(net25077), .B1(n343), .Y(n611));
sg13g2_nand2_2 U458 (.A(new_key_o_96_), .B(net25075), .Y(n343));
sg13g2_o21ai_1 U459 (.A1(n231), .A2(net25105), .B1(n232), .Y(n769));
sg13g2_o21ai_1 U460 (.A1(n345), .A2(net25107), .B1(n346), .Y(n612));
sg13g2_nand2_2 U461 (.A(new_key_o_128_), .B(net25075), .Y(n346));
sg13g2_inv_4 U462 (.A(n344), .Y(n345));
sg13g2_xnor2_1 U463 (.A(last_key_i_104_), .B(n810), .Y(n251));
sg13g2_o21ai_1 U464 (.A1(n347), .A2(net25127), .B1(n348), .Y(n613));
sg13g2_nand2_2 U465 (.A(new_key_o_160_), .B(net25075), .Y(n348));
sg13g2_o21ai_1 U466 (.A1(net25115), .A2(n74), .B1(n75), .Y(n717));
sg13g2_o21ai_1 U467 (.A1(net25111), .A2(n349), .B1(n350), .Y(n614));
sg13g2_nand2_2 U468 (.A(new_key_o_33_), .B(net25075), .Y(n350));
sg13g2_o21ai_1 U469 (.A1(n351), .A2(net25079), .B1(n352), .Y(n615));
sg13g2_nand2_2 U470 (.A(new_key_o_1_), .B(net25075), .Y(n352));
sg13g2_xnor2_1 U471 (.A(n39), .B(n349), .Y(n351));
sg13g2_xnor2_1 U472 (.A(n353), .B(last_key_i_33_), .Y(n349));
sg13g2_o21ai_1 U473 (.A1(n356), .A2(net25105), .B1(n357), .Y(n617));
sg13g2_o21ai_1 U474 (.A1(n354), .A2(net25103), .B1(n355), .Y(n616));
sg13g2_nand2_2 U475 (.A(new_key_o_65_), .B(net25075), .Y(n355));
sg13g2_inv_4 U476 (.A(n353), .Y(n354));
sg13g2_xnor2_1 U477 (.A(last_key_i_65_), .B(n356), .Y(n353));
sg13g2_xnor2_1 U478 (.A(last_key_i_97_), .B(n358), .Y(n356));
sg13g2_nand2_2 U479 (.A(new_key_o_97_), .B(net25075), .Y(n357));
sg13g2_inv_4 U480 (.A(n174), .Y(n175));
sg13g2_o21ai_1 U481 (.A1(n359), .A2(net25077), .B1(n360), .Y(n618));
sg13g2_nand2_2 U482 (.A(new_key_o_129_), .B(net25111), .Y(n360));
sg13g2_inv_4 U483 (.A(n358), .Y(n359));
sg13g2_o21ai_1 U484 (.A1(n169), .A2(net25115), .B1(n170), .Y(n746));
sg13g2_o21ai_1 U485 (.A1(n361), .A2(net25105), .B1(n362), .Y(n619));
sg13g2_nand2_2 U486 (.A(new_key_o_161_), .B(net25107), .Y(n362));
sg13g2_xnor2_1 U487 (.A(n344), .B(last_key_i_96_), .Y(n342));
sg13g2_xnor2_1 U488 (.A(n339), .B(last_key_i_32_), .Y(n335));
sg13g2_nand2_2 U489 (.A(new_key_o_34_), .B(net25105), .Y(n364));
sg13g2_xnor2_1 U490 (.A(last_key_i_64_), .B(n342), .Y(n339));
sg13g2_nand2_2 U491 (.A(new_key_o_2_), .B(net25109), .Y(n366));
sg13g2_inv_4 U492 (.A(last_key_i_61_), .Y(n963));
sg13g2_xnor2_1 U493 (.A(n497), .B(last_key_i_51_), .Y(n492));
sg13g2_o21ai_1 U494 (.A1(n477), .A2(net25113), .B1(n478), .Y(n668));
sg13g2_o21ai_1 U495 (.A1(net25081), .A2(n368), .B1(n369), .Y(n622));
sg13g2_nand2_2 U496 (.A(new_key_o_66_), .B(net25113), .Y(n369));
sg13g2_inv_4 U497 (.A(n367), .Y(n368));
sg13g2_xnor2_1 U498 (.A(n482), .B(last_key_i_50_), .Y(n477));
sg13g2_o21ai_1 U499 (.A1(n447), .A2(net25115), .B1(n448), .Y(n656));
sg13g2_nand2_2 U500 (.A(new_key_o_98_), .B(net25109), .Y(n371));
sg13g2_o21ai_1 U501 (.A1(n806), .A2(net25109), .B1(n525), .Y(n687));
sg13g2_o21ai_1 U502 (.A1(n373), .A2(net25107), .B1(n374), .Y(n624));
sg13g2_nand2_2 U503 (.A(new_key_o_130_), .B(net25111), .Y(n374));
sg13g2_nand2_2 U504 (.A(last_key_i_67_), .B(n384), .Y(n878));
sg13g2_o21ai_1 U505 (.A1(n384), .A2(net25081), .B1(n385), .Y(n629));
sg13g2_o21ai_1 U506 (.A1(net25115), .A2(n375), .B1(n376), .Y(n625));
sg13g2_nand2_2 U507 (.A(new_key_o_162_), .B(net25093), .Y(n376));
sg13g2_xnor2_1 U508 (.A(last_key_i_162_), .B(col_2), .Y(n375));
sg13g2_o21ai_1 U509 (.A1(n377), .A2(net25115), .B1(n378), .Y(n626));
sg13g2_nand2_2 U510 (.A(new_key_o_35_), .B(net25079), .Y(n378));
sg13g2_xnor2_1 U511 (.A(n386), .B(last_key_i_99_), .Y(n384));
sg13g2_nand2_2 U512 (.A(new_key_o_3_), .B(net25127), .Y(n380));
sg13g2_o21ai_1 U513 (.A1(n379), .A2(net25109), .B1(n380), .Y(n627));
sg13g2_xnor2_1 U514 (.A(n928), .B(n377), .Y(n379));
sg13g2_xnor2_1 U515 (.A(last_key_i_113_), .B(n472), .Y(n470));
sg13g2_o21ai_1 U516 (.A1(n382), .A2(net25093), .B1(n383), .Y(n628));
sg13g2_nand2_2 U517 (.A(new_key_o_67_), .B(net25075), .Y(n383));
sg13g2_inv_4 U518 (.A(n381), .Y(n382));
sg13g2_xnor2_1 U519 (.A(last_key_i_145_), .B(n475), .Y(n472));
sg13g2_inv_4 U520 (.A(last_key_i_0_), .Y(n44));
sg13g2_nand2_2 U521 (.A(new_key_o_99_), .B(net25093), .Y(n385));
sg13g2_inv_4 U522 (.A(last_key_i_6_), .Y(n14));
sg13g2_o21ai_1 U523 (.A1(n387), .A2(net25115), .B1(n388), .Y(n630));
sg13g2_nand2_2 U524 (.A(new_key_o_131_), .B(net25127), .Y(n388));
sg13g2_inv_4 U525 (.A(n386), .Y(n387));
sg13g2_inv_4 U526 (.A(last_key_i_4_), .Y(n24));
sg13g2_o21ai_1 U527 (.A1(n389), .A2(net25111), .B1(n390), .Y(n631));
sg13g2_nand2_2 U528 (.A(new_key_o_163_), .B(net25097), .Y(n390));
sg13g2_nand2_2 U529 (.A(n208), .B(last_key_i_41_), .Y(n812));
sg13g2_o21ai_1 U530 (.A1(n391), .A2(net25081), .B1(n392), .Y(n632));
sg13g2_nand2_2 U531 (.A(new_key_o_36_), .B(net25083), .Y(n392));
sg13g2_nand2_2 U532 (.A(n206), .B(n811), .Y(n813));
sg13g2_nand2_2 U533 (.A(new_key_o_4_), .B(net25127), .Y(n394));
sg13g2_nand2_2 U534 (.A(n813), .B(n812), .Y(n224));
sg13g2_inv_4 U535 (.A(last_key_i_41_), .Y(n811));
sg13g2_inv_4 U536 (.A(n196), .Y(n194));
sg13g2_o21ai_1 U537 (.A1(n396), .A2(net25109), .B1(n397), .Y(n634));
sg13g2_nand2_2 U538 (.A(new_key_o_68_), .B(net25081), .Y(n397));
sg13g2_inv_4 U539 (.A(n395), .Y(n396));
sg13g2_xnor2_1 U540 (.A(last_key_i_31_), .B(n169), .Y(n173));
sg13g2_o21ai_1 U541 (.A1(n398), .A2(net25075), .B1(n399), .Y(n635));
sg13g2_nand2_2 U542 (.A(new_key_o_100_), .B(net25113), .Y(n399));
sg13g2_nand2_2 U543 (.A(sbox_data_i_3_), .B(last_key_i_171_), .Y(n899));
sg13g2_o21ai_1 U544 (.A1(n401), .A2(net25113), .B1(n402), .Y(n636));
sg13g2_nand2_2 U545 (.A(new_key_o_132_), .B(net25093), .Y(n402));
sg13g2_inv_4 U546 (.A(n400), .Y(n401));
sg13g2_nand2_2 U547 (.A(n226), .B(n984), .Y(n815));
sg13g2_o21ai_1 U548 (.A1(n403), .A2(net25079), .B1(n404), .Y(n637));
sg13g2_nand2_2 U549 (.A(new_key_o_164_), .B(net25077), .Y(n404));
sg13g2_nand2_2 U550 (.A(n814), .B(last_key_i_8_), .Y(n816));
sg13g2_o21ai_1 U551 (.A1(n405), .A2(net25103), .B1(n406), .Y(n638));
sg13g2_nand2_2 U552 (.A(new_key_o_37_), .B(net25107), .Y(n406));
sg13g2_o21ai_1 U553 (.A1(n407), .A2(net25107), .B1(n408), .Y(n639));
sg13g2_nand2_2 U554 (.A(new_key_o_5_), .B(net25107), .Y(n408));
sg13g2_xnor2_1 U555 (.A(n19), .B(n405), .Y(n407));
sg13g2_nand2_2 U556 (.A(n815), .B(n816), .Y(n249));
sg13g2_inv_4 U557 (.A(n226), .Y(n814));
sg13g2_o21ai_1 U558 (.A1(n410), .A2(net25127), .B1(n411), .Y(n640));
sg13g2_nand2_2 U559 (.A(new_key_o_69_), .B(net25079), .Y(n411));
sg13g2_inv_4 U560 (.A(n409), .Y(n410));
sg13g2_inv_4 U561 (.A(round_i_3_), .Y(n187));
sg13g2_o21ai_1 U562 (.A1(n412), .A2(net25105), .B1(n413), .Y(n641));
sg13g2_nand2_2 U563 (.A(new_key_o_101_), .B(net25081), .Y(n413));
sg13g2_nand2_2 U564 (.A(sbox_data_i_2_), .B(last_key_i_170_), .Y(n820));
sg13g2_o21ai_1 U565 (.A1(n415), .A2(net25075), .B1(n416), .Y(n642));
sg13g2_nand2_2 U566 (.A(new_key_o_133_), .B(net25083), .Y(n416));
sg13g2_inv_4 U567 (.A(n904), .Y(n415));
sg13g2_nand2_2 U568 (.A(n818), .B(n819), .Y(n821));
sg13g2_o21ai_1 U569 (.A1(n417), .A2(net25115), .B1(n418), .Y(n643));
sg13g2_nand2_2 U570 (.A(new_key_o_165_), .B(net25103), .Y(n418));
sg13g2_nand2_2 U571 (.A(n820), .B(n821), .Y(n276));
sg13g2_inv_4 U572 (.A(last_key_i_170_), .Y(n818));
sg13g2_nand2_2 U573 (.A(new_key_o_38_), .B(net25111), .Y(n420));
sg13g2_o21ai_1 U574 (.A1(n421), .A2(net25103), .B1(n422), .Y(n645));
sg13g2_nand2_2 U575 (.A(new_key_o_6_), .B(net25075), .Y(n422));
sg13g2_xnor2_1 U576 (.A(n14), .B(n419), .Y(n421));
sg13g2_inv_4 U577 (.A(sbox_data_i_2_), .Y(n819));
sg13g2_o21ai_1 U578 (.A1(n249), .A2(net25127), .B1(n250), .Y(n775));
sg13g2_o21ai_1 U579 (.A1(n874), .A2(net25111), .B1(n425), .Y(n646));
sg13g2_nand2_2 U580 (.A(new_key_o_70_), .B(net25079), .Y(n425));
sg13g2_nand2_2 U581 (.A(n899), .B(n808), .Y(n822));
sg13g2_xnor2_1 U582 (.A(n214), .B(n10), .Y(n231));
sg13g2_nand2_2 U583 (.A(n224), .B(n35), .Y(n824));
sg13g2_nand2_2 U584 (.A(new_key_o_102_), .B(net25113), .Y(n427));
sg13g2_nand2_2 U585 (.A(n823), .B(n839), .Y(n825));
sg13g2_o21ai_1 U586 (.A1(n429), .A2(net25113), .B1(n430), .Y(n648));
sg13g2_nand2_2 U587 (.A(new_key_o_134_), .B(net25103), .Y(n430));
sg13g2_inv_4 U588 (.A(n428), .Y(n429));
sg13g2_nand2_2 U589 (.A(n825), .B(n824), .Y(n246));
sg13g2_o21ai_1 U590 (.A1(n431), .A2(net25097), .B1(n432), .Y(n649));
sg13g2_nand2_2 U591 (.A(new_key_o_166_), .B(net25097), .Y(n432));
sg13g2_inv_4 U592 (.A(n224), .Y(n823));
sg13g2_nand3_1 U593 (.A(n11), .B(n990), .C(n12), .Y(sbox_data_o_6_));
sg13g2_nand2_2 U594 (.A(new_key_o_39_), .B(net25097), .Y(n434));
sg13g2_inv_4 U595 (.A(last_key_i_14_), .Y(n10));
sg13g2_nand2_2 U596 (.A(new_key_o_7_), .B(net25127), .Y(n436));
sg13g2_xnor2_1 U597 (.A(last_key_i_142_), .B(n288), .Y(n265));
sg13g2_nand2_2 U598 (.A(sbox_data_i_4_), .B(last_key_i_172_), .Y(n829));
sg13g2_nand2_2 U599 (.A(n827), .B(n828), .Y(n830));
sg13g2_o21ai_1 U600 (.A1(net25115), .A2(n438), .B1(n439), .Y(n652));
sg13g2_nand2_2 U601 (.A(new_key_o_71_), .B(net25093), .Y(n439));
sg13g2_inv_4 U602 (.A(n437), .Y(n438));
sg13g2_xnor2_1 U603 (.A(n440), .B(last_key_i_71_), .Y(n437));
sg13g2_o21ai_1 U604 (.A1(net25115), .A2(n440), .B1(n441), .Y(n653));
sg13g2_nand2_2 U605 (.A(new_key_o_103_), .B(net25107), .Y(n441));
sg13g2_nand2_2 U606 (.A(n829), .B(n830), .Y(n282));
sg13g2_o21ai_1 U607 (.A1(n443), .A2(net25115), .B1(n444), .Y(n654));
sg13g2_nand2_2 U608 (.A(new_key_o_135_), .B(net25111), .Y(n444));
sg13g2_inv_4 U609 (.A(n442), .Y(n443));
sg13g2_xnor2_1 U610 (.A(n233), .B(last_key_i_78_), .Y(n193));
sg13g2_o21ai_1 U611 (.A1(net25115), .A2(n445), .B1(n446), .Y(n655));
sg13g2_nand2_2 U612 (.A(new_key_o_167_), .B(net25097), .Y(n446));
sg13g2_nand2_2 U613 (.A(n236), .B(last_key_i_77_), .Y(n833));
sg13g2_nand2_2 U614 (.A(n832), .B(n831), .Y(n834));
sg13g2_nand2_2 U615 (.A(new_key_o_48_), .B(net25103), .Y(n448));
sg13g2_nand2_2 U616 (.A(n833), .B(n834), .Y(n196));
sg13g2_nand2_2 U617 (.A(new_key_o_16_), .B(net25097), .Y(n450));
sg13g2_inv_4 U618 (.A(n451), .Y(n449));
sg13g2_xnor2_1 U619 (.A(last_key_i_16_), .B(n447), .Y(n451));
sg13g2_inv_4 U620 (.A(last_key_i_77_), .Y(n831));
sg13g2_o21ai_1 U621 (.A1(n453), .A2(net25115), .B1(n454), .Y(n658));
sg13g2_nand2_2 U622 (.A(new_key_o_80_), .B(net25109), .Y(n454));
sg13g2_inv_4 U623 (.A(n452), .Y(n453));
sg13g2_inv_4 U624 (.A(n236), .Y(n832));
sg13g2_o21ai_1 U625 (.A1(n455), .A2(net25115), .B1(n456), .Y(n659));
sg13g2_nand2_2 U626 (.A(new_key_o_112_), .B(net25079), .Y(n456));
sg13g2_o21ai_1 U627 (.A1(n214), .A2(net25103), .B1(n215), .Y(n761));
sg13g2_o21ai_1 U628 (.A1(n458), .A2(net25115), .B1(n459), .Y(n660));
sg13g2_nand2_2 U629 (.A(new_key_o_144_), .B(net25075), .Y(n459));
sg13g2_inv_4 U630 (.A(n457), .Y(n458));
sg13g2_nand2_2 U631 (.A(last_key_i_74_), .B(n245), .Y(n837));
sg13g2_o21ai_1 U632 (.A1(n804), .A2(net25115), .B1(n461), .Y(n661));
sg13g2_nand2_2 U633 (.A(new_key_o_176_), .B(net25097), .Y(n461));
sg13g2_nand2_2 U634 (.A(n837), .B(n838), .Y(n205));
sg13g2_o21ai_1 U635 (.A1(n462), .A2(net25113), .B1(n463), .Y(n662));
sg13g2_nand2_2 U636 (.A(new_key_o_49_), .B(net25113), .Y(n463));
sg13g2_inv_4 U637 (.A(n245), .Y(n836));
sg13g2_nand2_2 U638 (.A(new_key_o_17_), .B(net25115), .Y(n465));
sg13g2_inv_4 U639 (.A(n466), .Y(n464));
sg13g2_xnor2_1 U640 (.A(last_key_i_17_), .B(n462), .Y(n466));
sg13g2_xnor2_1 U641 (.A(last_key_i_42_), .B(n205), .Y(n222));
sg13g2_o21ai_1 U642 (.A1(n468), .A2(net25113), .B1(n469), .Y(n664));
sg13g2_nand2_2 U643 (.A(new_key_o_81_), .B(net25097), .Y(n469));
sg13g2_inv_4 U644 (.A(n467), .Y(n468));
sg13g2_inv_4 U645 (.A(n35), .Y(n839));
sg13g2_o21ai_1 U646 (.A1(n470), .A2(net25113), .B1(n471), .Y(n665));
sg13g2_nand2_2 U647 (.A(new_key_o_113_), .B(net25127), .Y(n471));
sg13g2_inv_4 U648 (.A(last_key_i_9_), .Y(n35));
sg13g2_o21ai_1 U649 (.A1(n473), .A2(net25113), .B1(n474), .Y(n666));
sg13g2_nand2_2 U650 (.A(new_key_o_145_), .B(net25097), .Y(n474));
sg13g2_inv_4 U651 (.A(n472), .Y(n473));
sg13g2_nand2_2 U652 (.A(n196), .B(last_key_i_45_), .Y(n841));
sg13g2_o21ai_1 U653 (.A1(n475), .A2(net25113), .B1(n476), .Y(n667));
sg13g2_nand2_2 U654 (.A(new_key_o_177_), .B(net25081), .Y(n476));
sg13g2_nand2_2 U655 (.A(n194), .B(n840), .Y(n842));
sg13g2_nand2_2 U656 (.A(n842), .B(n841), .Y(n216));
sg13g2_nand2_2 U657 (.A(new_key_o_50_), .B(net25097), .Y(n478));
sg13g2_o21ai_1 U658 (.A1(n479), .A2(net25113), .B1(n480), .Y(n669));
sg13g2_nand2_2 U659 (.A(new_key_o_18_), .B(net25113), .Y(n480));
sg13g2_inv_4 U660 (.A(last_key_i_45_), .Y(n840));
sg13g2_nand2_2 U661 (.A(n844), .B(n843), .Y(n846));
sg13g2_inv_4 U662 (.A(last_key_i_136_), .Y(n843));
sg13g2_o21ai_1 U663 (.A1(n483), .A2(net25113), .B1(n484), .Y(n670));
sg13g2_nand2_2 U664 (.A(new_key_o_82_), .B(net25083), .Y(n484));
sg13g2_inv_4 U665 (.A(n482), .Y(n483));
sg13g2_inv_4 U666 (.A(n817), .Y(n844));
sg13g2_o21ai_1 U667 (.A1(n485), .A2(net25113), .B1(n486), .Y(n671));
sg13g2_nand2_2 U668 (.A(new_key_o_114_), .B(net25097), .Y(n486));
sg13g2_nand2_2 U669 (.A(n251), .B(last_key_i_72_), .Y(n849));
sg13g2_o21ai_1 U670 (.A1(n914), .A2(net25113), .B1(n489), .Y(n672));
sg13g2_nand2_2 U671 (.A(new_key_o_146_), .B(net25081), .Y(n489));
sg13g2_nand2_2 U672 (.A(n848), .B(n847), .Y(n850));
sg13g2_nand2_2 U673 (.A(n849), .B(n850), .Y(n211));
sg13g2_o21ai_1 U674 (.A1(n490), .A2(net25113), .B1(n491), .Y(n673));
sg13g2_nand2_2 U675 (.A(new_key_o_178_), .B(net25093), .Y(n491));
sg13g2_xnor2_1 U676 (.A(last_key_i_178_), .B(col_18_), .Y(n490));
sg13g2_o21ai_1 U677 (.A1(n492), .A2(net25111), .B1(n493), .Y(n674));
sg13g2_nand2_2 U678 (.A(new_key_o_51_), .B(net25093), .Y(n493));
sg13g2_inv_4 U679 (.A(last_key_i_72_), .Y(n847));
sg13g2_nand2_2 U680 (.A(new_key_o_19_), .B(net25093), .Y(n495));
sg13g2_inv_4 U681 (.A(n251), .Y(n848));
sg13g2_o21ai_1 U682 (.A1(n237), .A2(net25105), .B1(n238), .Y(n771));
sg13g2_o21ai_1 U683 (.A1(n240), .A2(net25105), .B1(n241), .Y(n772));
sg13g2_o21ai_1 U684 (.A1(n498), .A2(net25111), .B1(n499), .Y(n676));
sg13g2_nand2_2 U685 (.A(new_key_o_83_), .B(net25093), .Y(n499));
sg13g2_inv_4 U686 (.A(n497), .Y(n498));
sg13g2_xnor2_1 U687 (.A(n174), .B(last_key_i_63_), .Y(n169));
sg13g2_o21ai_1 U688 (.A1(n500), .A2(net25111), .B1(n501), .Y(n677));
sg13g2_nand2_2 U689 (.A(new_key_o_115_), .B(net25093), .Y(n501));
sg13g2_xnor2_1 U690 (.A(last_key_i_43_), .B(n202), .Y(n220));
sg13g2_o21ai_1 U691 (.A1(n907), .A2(net25111), .B1(n504), .Y(n678));
sg13g2_nand2_2 U692 (.A(new_key_o_147_), .B(net25093), .Y(n504));
sg13g2_nand3_1 U693 (.A(n50), .B(n318), .C(n49), .Y(n301));
sg13g2_inv_4 U694 (.A(n248), .Y(n981));
sg13g2_o21ai_1 U695 (.A1(n505), .A2(net25111), .B1(n506), .Y(n679));
sg13g2_nand2_2 U696 (.A(new_key_o_179_), .B(net25083), .Y(n506));
sg13g2_o21ai_1 U697 (.A1(n822), .A2(net25109), .B1(n295), .Y(n795));
sg13g2_o21ai_1 U698 (.A1(n507), .A2(net25111), .B1(n508), .Y(n680));
sg13g2_nand2_2 U699 (.A(new_key_o_52_), .B(net25077), .Y(n508));
sg13g2_o21ai_1 U700 (.A1(n509), .A2(net25111), .B1(n510), .Y(n681));
sg13g2_nand2_2 U701 (.A(new_key_o_20_), .B(net25111), .Y(n510));
sg13g2_inv_4 U702 (.A(n511), .Y(n509));
sg13g2_xnor2_1 U703 (.A(last_key_i_20_), .B(n507), .Y(n511));
sg13g2_o21ai_1 U704 (.A1(net25113), .A2(n312), .B1(n297), .Y(n797));
sg13g2_o21ai_1 U705 (.A1(n513), .A2(net25111), .B1(n514), .Y(n682));
sg13g2_nand2_2 U706 (.A(new_key_o_84_), .B(net25081), .Y(n514));
sg13g2_inv_4 U707 (.A(n512), .Y(n513));
sg13g2_nand2_2 U708 (.A(last_key_i_23_), .B(n9), .Y(n3));
sg13g2_o21ai_1 U709 (.A1(n515), .A2(net25111), .B1(n516), .Y(n683));
sg13g2_nand2_2 U710 (.A(new_key_o_116_), .B(net25107), .Y(n516));
sg13g2_inv_4 U711 (.A(n7), .Y(n855));
sg13g2_o21ai_1 U712 (.A1(n936), .A2(net25111), .B1(n519), .Y(n684));
sg13g2_nand2_2 U713 (.A(new_key_o_148_), .B(net25083), .Y(n519));
sg13g2_nor2_2 U714 (.A(n34), .B(n7), .Y(n33));
sg13g2_nand3_1 U715 (.A(state_0_), .B(n318), .C(state_1_), .Y(n7));
sg13g2_o21ai_1 U716 (.A1(n520), .A2(net25111), .B1(n521), .Y(n685));
sg13g2_nand2_2 U717 (.A(new_key_o_180_), .B(net25111), .Y(n521));
sg13g2_nand2_2 U718 (.A(last_key_i_16_), .B(n9), .Y(n41));
sg13g2_o21ai_1 U719 (.A1(n522), .A2(net25109), .B1(n523), .Y(n686));
sg13g2_nand2_2 U720 (.A(new_key_o_53_), .B(net25077), .Y(n523));
sg13g2_nand2_2 U721 (.A(n248), .B(last_key_i_73_), .Y(n982));
sg13g2_nand2_2 U722 (.A(new_key_o_21_), .B(net25081), .Y(n525));
sg13g2_nand2_2 U723 (.A(n981), .B(n980), .Y(n983));
sg13g2_o21ai_1 U724 (.A1(n218), .A2(n943), .B1(n888), .Y(n237));
sg13g2_nand4_1 U725 (.A(n47), .B(net39263), .C(n48), .D(n7), .Y(sbox_access_o));
sg13g2_o21ai_1 U726 (.A1(n929), .A2(net25109), .B1(n529), .Y(n688));
sg13g2_nand2_2 U727 (.A(new_key_o_85_), .B(net25081), .Y(n529));
sg13g2_nand2_2 U728 (.A(last_key_i_4_), .B(n855), .Y(n856));
sg13g2_inv_4 U729 (.A(n45), .Y(n9));
sg13g2_o21ai_1 U730 (.A1(net25109), .A2(n530), .B1(n531), .Y(n689));
sg13g2_nand2_2 U731 (.A(new_key_o_117_), .B(net25075), .Y(n531));
sg13g2_nand2_2 U732 (.A(last_key_i_6_), .B(n855), .Y(n857));
sg13g2_o21ai_1 U733 (.A1(n533), .A2(net25109), .B1(n534), .Y(n690));
sg13g2_nand2_2 U734 (.A(new_key_o_149_), .B(net25127), .Y(n534));
sg13g2_inv_4 U735 (.A(n532), .Y(n533));
sg13g2_inv_4 U736 (.A(n857), .Y(n13));
sg13g2_o21ai_1 U737 (.A1(n535), .A2(net25109), .B1(n536), .Y(n691));
sg13g2_nand2_2 U738 (.A(new_key_o_181_), .B(net25097), .Y(n536));
sg13g2_nand3_1 U739 (.A(n31), .B(n991), .C(n32), .Y(sbox_data_o_2_));
sg13g2_o21ai_1 U740 (.A1(n537), .A2(net25109), .B1(n538), .Y(n692));
sg13g2_nand2_2 U741 (.A(new_key_o_54_), .B(net25127), .Y(n538));
sg13g2_nor2_2 U742 (.A(n300), .B(n301), .Y(n5));
sg13g2_nand2_2 U743 (.A(new_key_o_22_), .B(net25083), .Y(n540));
sg13g2_inv_4 U744 (.A(last_key_i_30_), .Y(net25830));
sg13g2_nand2_2 U745 (.A(last_key_i_22_), .B(n9), .Y(n11));
sg13g2_inv_4 U746 (.A(last_key_i_26_), .Y(n858));
sg13g2_o21ai_1 U747 (.A1(n543), .A2(net25109), .B1(n544), .Y(n694));
sg13g2_nand2_2 U748 (.A(new_key_o_86_), .B(net25097), .Y(n544));
sg13g2_inv_4 U749 (.A(n542), .Y(n543));
sg13g2_inv_4 U750 (.A(n858), .Y(n859));
sg13g2_inv_4 U751 (.A(last_key_i_7_), .Y(n8));
sg13g2_nand2_2 U752 (.A(new_key_o_118_), .B(net25107), .Y(n546));
sg13g2_xnor2_1 U753 (.A(last_key_i_188_), .B(col_28_), .Y(n129));
sg13g2_o21ai_1 U754 (.A1(n548), .A2(net25109), .B1(n549), .Y(n696));
sg13g2_nand2_2 U755 (.A(new_key_o_150_), .B(net25093), .Y(n549));
sg13g2_inv_4 U756 (.A(n547), .Y(n548));
sg13g2_xnor2_1 U757 (.A(n550), .B(last_key_i_150_), .Y(n547));
sg13g2_o21ai_1 U758 (.A1(net25109), .A2(n550), .B1(n551), .Y(n697));
sg13g2_nand2_2 U759 (.A(new_key_o_182_), .B(net25075), .Y(n551));
sg13g2_xnor2_1 U760 (.A(last_key_i_182_), .B(col_22_), .Y(n550));
sg13g2_o21ai_1 U761 (.A1(n552), .A2(net25107), .B1(n553), .Y(n698));
sg13g2_nand2_2 U762 (.A(new_key_o_55_), .B(net25081), .Y(n553));
sg13g2_nand2_2 U763 (.A(last_key_i_87_), .B(n560), .Y(n860));
sg13g2_nand2_2 U764 (.A(new_key_o_23_), .B(net25077), .Y(n555));
sg13g2_nand2_2 U765 (.A(n562), .B(last_key_i_119_), .Y(n862));
sg13g2_nand2_2 U766 (.A(n563), .B(n861), .Y(n863));
sg13g2_nand2_2 U767 (.A(n862), .B(n863), .Y(n560));
sg13g2_o21ai_1 U768 (.A1(n558), .A2(net25107), .B1(n559), .Y(n700));
sg13g2_nand2_2 U769 (.A(new_key_o_87_), .B(net25077), .Y(n559));
sg13g2_inv_4 U770 (.A(n557), .Y(n558));
sg13g2_inv_4 U771 (.A(last_key_i_119_), .Y(n861));
sg13g2_xnor2_1 U772 (.A(n557), .B(last_key_i_55_), .Y(n552));
sg13g2_nand2_2 U773 (.A(new_key_o_119_), .B(net25111), .Y(n561));
sg13g2_o21ai_1 U774 (.A1(n560), .A2(net25107), .B1(n561), .Y(n701));
sg13g2_o21ai_1 U775 (.A1(n563), .A2(net25107), .B1(n564), .Y(n702));
sg13g2_nand2_2 U776 (.A(new_key_o_151_), .B(net25113), .Y(n564));
sg13g2_xnor2_1 U777 (.A(last_key_i_68_), .B(n398), .Y(n395));
sg13g2_xnor2_1 U778 (.A(last_key_i_100_), .B(n400), .Y(n398));
sg13g2_o21ai_1 U779 (.A1(n565), .A2(net25107), .B1(n566), .Y(n703));
sg13g2_nand2_2 U780 (.A(new_key_o_183_), .B(net25077), .Y(n566));
sg13g2_xnor2_1 U781 (.A(last_key_i_69_), .B(n412), .Y(n409));
sg13g2_o21ai_1 U782 (.A1(n567), .A2(net25107), .B1(n568), .Y(n704));
sg13g2_nand2_2 U783 (.A(new_key_o_56_), .B(net25075), .Y(n568));
sg13g2_xnor2_1 U784 (.A(last_key_i_101_), .B(n904), .Y(n412));
sg13g2_nand2_2 U785 (.A(new_key_o_24_), .B(net25097), .Y(n570));
sg13g2_nand3_1 U786 (.A(n89), .B(n110), .C(n150), .Y(n148));
sg13g2_nand4_1 U787 (.A(n130), .B(n109), .C(n89), .D(n70), .Y(n128));
sg13g2_nand2_2 U788 (.A(n437), .B(last_key_i_39_), .Y(n869));
sg13g2_o21ai_1 U789 (.A1(n573), .A2(net25107), .B1(n574), .Y(n706));
sg13g2_nand2_2 U790 (.A(new_key_o_88_), .B(net25083), .Y(n574));
sg13g2_inv_4 U791 (.A(n572), .Y(n573));
sg13g2_nand2_2 U792 (.A(n869), .B(n870), .Y(n433));
sg13g2_o21ai_1 U793 (.A1(n575), .A2(net25107), .B1(n576), .Y(n707));
sg13g2_nand2_2 U794 (.A(new_key_o_120_), .B(net25081), .Y(n576));
sg13g2_inv_4 U795 (.A(last_key_i_39_), .Y(n868));
sg13g2_o21ai_1 U796 (.A1(n578), .A2(net25077), .B1(n579), .Y(n708));
sg13g2_nand2_2 U797 (.A(new_key_o_152_), .B(net25083), .Y(n579));
sg13g2_inv_4 U798 (.A(n577), .Y(n578));
sg13g2_o21ai_1 U799 (.A1(n435), .A2(net25115), .B1(n436), .Y(n651));
sg13g2_o21ai_1 U800 (.A1(n580), .A2(net25107), .B1(n581), .Y(n709));
sg13g2_nand2_2 U801 (.A(new_key_o_184_), .B(net25093), .Y(n581));
sg13g2_nand3_1 U802 (.A(n49), .B(n50), .C(n301), .Y(n52));
sg13g2_o21ai_1 U803 (.A1(n433), .A2(net25115), .B1(n434), .Y(n650));
sg13g2_a21oi_1 U804 (.A1(n992), .A2(n88), .B1(n186), .Y(n184));
sg13g2_nand2_2 U805 (.A(n428), .B(last_key_i_102_), .Y(n872));
sg13g2_nand2_2 U806 (.A(n872), .B(n873), .Y(n426));
sg13g2_inv_4 U807 (.A(last_key_i_102_), .Y(n871));
sg13g2_nand2_2 U808 (.A(n90), .B(n132), .Y(n582));
sg13g2_nand2_2 U809 (.A(n423), .B(last_key_i_38_), .Y(n876));
sg13g2_nand2_2 U810 (.A(n874), .B(n875), .Y(n877));
sg13g2_nand2_2 U811 (.A(n876), .B(n877), .Y(n419));
sg13g2_inv_4 U812 (.A(n423), .Y(n874));
sg13g2_inv_4 U813 (.A(last_key_i_38_), .Y(n875));
sg13g2_xnor2_1 U814 (.A(last_key_i_70_), .B(n426), .Y(n423));
sg13g2_o21ai_1 U815 (.A1(n426), .A2(net25105), .B1(n427), .Y(n647));
sg13g2_o21ai_1 U816 (.A1(n419), .A2(net25115), .B1(n420), .Y(n644));
sg13g2_nand2_2 U817 (.A(last_key_i_163_), .B(col_3), .Y(n881));
sg13g2_nand2_2 U818 (.A(n879), .B(n880), .Y(n882));
sg13g2_nand2_2 U819 (.A(n881), .B(n882), .Y(n389));
sg13g2_inv_4 U820 (.A(last_key_i_163_), .Y(n879));
sg13g2_and2_1 U821 (.A(n111), .B(n131), .X(n992));
sg13g2_xnor2_1 U822 (.A(n381), .B(last_key_i_35_), .Y(n377));
sg13g2_nand2_2 U823 (.A(n34), .B(n363), .Y(n885));
sg13g2_nand2_2 U824 (.A(n883), .B(n884), .Y(n886));
sg13g2_nand2_2 U825 (.A(n886), .B(n885), .Y(n365));
sg13g2_inv_4 U826 (.A(n34), .Y(n883));
sg13g2_inv_4 U827 (.A(n363), .Y(n884));
sg13g2_nand2_2 U828 (.A(n367), .B(last_key_i_34_), .Y(n887));
sg13g2_inv_4 U829 (.A(last_key_i_2_), .Y(n34));
sg13g2_o21ai_1 U830 (.A1(n365), .A2(net25077), .B1(n366), .Y(n621));
sg13g2_o21ai_1 U831 (.A1(n363), .A2(net25097), .B1(n364), .Y(n620));
sg13g2_xnor2_1 U832 (.A(last_key_i_160_), .B(col_0), .Y(n347));
sg13g2_o21ai_1 U833 (.A1(n69), .A2(n88), .B1(n89), .Y(n86));
sg13g2_nand2_2 U834 (.A(round_i_1_), .B(n90), .Y(n69));
sg13g2_nand2_2 U835 (.A(sbox_data_i_5_), .B(last_key_i_173_), .Y(n891));
sg13g2_nand2_2 U836 (.A(n889), .B(n890), .Y(n892));
sg13g2_inv_4 U837 (.A(sbox_data_i_5_), .Y(n889));
sg13g2_inv_1 U838 (.A(n1), .Y(n993));
sg13g2_nor2_2 U839 (.A(n88), .B(round_i_1_), .Y(n132));
sg13g2_inv_4 U840 (.A(last_key_i_13_), .Y(n15));
sg13g2_inv_4 U841 (.A(last_key_i_5_), .Y(n19));
sg13g2_nand4_1 U842 (.A(n108), .B(n109), .C(n70), .D(n110), .Y(n106));
sg13g2_o21ai_1 U843 (.A1(net25109), .A2(n94), .B1(n95), .Y(n723));
sg13g2_xnor2_1 U844 (.A(n957), .B(n93), .Y(n94));
sg13g2_nand2_2 U845 (.A(n242), .B(last_key_i_75_), .Y(n895));
sg13g2_nand2_2 U846 (.A(n894), .B(n893), .Y(n896));
sg13g2_nand2_2 U847 (.A(n895), .B(n896), .Y(n202));
sg13g2_inv_4 U848 (.A(n242), .Y(n894));
sg13g2_nand2_2 U849 (.A(n808), .B(n899), .Y(n279));
sg13g2_xnor2_1 U850 (.A(last_key_i_180_), .B(col_20_), .Y(n520));
sg13g2_nand2_2 U851 (.A(last_key_i_148_), .B(n520), .Y(n941));
sg13g2_xnor2_1 U852 (.A(last_key_i_52_), .B(n512), .Y(n507));
sg13g2_nand2_2 U853 (.A(last_key_i_86_), .B(n545), .Y(n900));
sg13g2_nand2_2 U854 (.A(n547), .B(last_key_i_118_), .Y(n902));
sg13g2_nand2_2 U855 (.A(n548), .B(n901), .Y(n903));
sg13g2_nand2_2 U856 (.A(n902), .B(n903), .Y(n545));
sg13g2_inv_4 U857 (.A(last_key_i_118_), .Y(n901));
sg13g2_xnor2_1 U858 (.A(n542), .B(last_key_i_54_), .Y(n537));
sg13g2_o21ai_1 U859 (.A1(n545), .A2(net25109), .B1(n546), .Y(n695));
sg13g2_nand2_1 U860 (.A(last_key_i_15_), .B(n993), .Y(n988));
sg13g2_a21oi_2 U861 (.A1(last_key_i_31_), .A2(net39266), .B1(n6), .Y(n4));
sg13g2_nor2_2 U862 (.A(n8), .B(n7), .Y(n6));
sg13g2_inv_4 U863 (.A(n8), .Y(net26231));
sg13g2_inv_4 U864 (.A(last_key_i_15_), .Y(n2));
sg13g2_inv_4 U865 (.A(last_key_i_23_), .Y(net25888));
sg13g2_xnor2_1 U866 (.A(last_key_i_165_), .B(col_5), .Y(n417));
sg13g2_xnor2_1 U867 (.A(last_key_i_129_), .B(n361), .Y(n358));
sg13g2_xnor2_1 U868 (.A(last_key_i_161_), .B(col_1), .Y(n361));
sg13g2_inv_4 U869 (.A(last_key_i_19_), .Y(n905));
sg13g2_inv_4 U870 (.A(n905), .Y(n906));
sg13g2_a21oi_2 U871 (.A1(last_key_i_27_), .A2(net39266), .B1(n28), .Y(n27));
sg13g2_nor2_2 U872 (.A(n29), .B(n7), .Y(n28));
sg13g2_nand2_2 U873 (.A(last_key_i_115_), .B(n502), .Y(n908));
sg13g2_nand2_2 U874 (.A(last_key_i_147_), .B(n505), .Y(n911));
sg13g2_nand2_2 U875 (.A(n909), .B(n910), .Y(n912));
sg13g2_nand2_2 U876 (.A(n911), .B(n912), .Y(n502));
sg13g2_inv_4 U877 (.A(last_key_i_147_), .Y(n909));
sg13g2_inv_4 U878 (.A(n505), .Y(n910));
sg13g2_xnor2_1 U879 (.A(last_key_i_83_), .B(n500), .Y(n497));
sg13g2_nand2_2 U880 (.A(last_key_i_114_), .B(n487), .Y(n915));
sg13g2_nand2_2 U881 (.A(n915), .B(n916), .Y(n485));
sg13g2_inv_4 U882 (.A(last_key_i_114_), .Y(n913));
sg13g2_nand2_2 U883 (.A(last_key_i_146_), .B(n490), .Y(n919));
sg13g2_nand2_2 U884 (.A(n919), .B(n920), .Y(n487));
sg13g2_inv_4 U885 (.A(last_key_i_146_), .Y(n917));
sg13g2_inv_4 U886 (.A(n490), .Y(n918));
sg13g2_xnor2_1 U887 (.A(last_key_i_82_), .B(n485), .Y(n482));
sg13g2_o21ai_1 U888 (.A1(net25105), .A2(n136), .B1(n137), .Y(n735));
sg13g2_o21ai_1 U889 (.A1(n464), .A2(net25113), .B1(n465), .Y(n663));
sg13g2_o21ai_1 U890 (.A1(net25111), .A2(n171), .B1(n172), .Y(n747));
sg13g2_nand2_2 U891 (.A(last_key_i_112_), .B(n457), .Y(n921));
sg13g2_nand2_2 U892 (.A(last_key_i_144_), .B(n804), .Y(n924));
sg13g2_nand2_2 U893 (.A(n922), .B(n923), .Y(n925));
sg13g2_nand2_2 U894 (.A(n924), .B(n925), .Y(n457));
sg13g2_inv_4 U895 (.A(last_key_i_144_), .Y(n922));
sg13g2_xnor2_1 U896 (.A(last_key_i_80_), .B(n455), .Y(n452));
sg13g2_xnor2_1 U897 (.A(last_key_i_139_), .B(n279), .Y(n259));
sg13g2_xnor2_1 U898 (.A(last_key_i_137_), .B(n273), .Y(n255));
sg13g2_xnor2_1 U899 (.A(last_key_i_138_), .B(n276), .Y(n257));
sg13g2_o21ai_1 U900 (.A1(n246), .A2(net25127), .B1(n247), .Y(n774));
sg13g2_xnor2_1 U901 (.A(last_key_i_56_), .B(n572), .Y(n567));
sg13g2_xnor2_1 U902 (.A(last_key_i_88_), .B(n575), .Y(n572));
sg13g2_inv_4 U903 (.A(last_key_i_21_), .Y(n926));
sg13g2_inv_4 U904 (.A(n29), .Y(n927));
sg13g2_inv_4 U905 (.A(n927), .Y(n928));
sg13g2_xnor2_1 U906 (.A(col_31_), .B(last_key_i_191_), .Y(n185));
sg13g2_a21oi_2 U907 (.A1(last_key_i_26_), .A2(net39266), .B1(n33), .Y(n32));
sg13g2_xnor2_1 U908 (.A(n184), .B(n185), .Y(n182));
sg13g2_nand2_2 U909 (.A(last_key_i_53_), .B(n527), .Y(n930));
sg13g2_nand2_2 U910 (.A(last_key_i_85_), .B(n530), .Y(n933));
sg13g2_nand2_2 U911 (.A(n933), .B(n934), .Y(n527));
sg13g2_inv_4 U912 (.A(last_key_i_85_), .Y(n931));
sg13g2_inv_4 U913 (.A(n530), .Y(n932));
sg13g2_nand2_2 U914 (.A(last_key_i_116_), .B(n517), .Y(n937));
sg13g2_nand2_2 U915 (.A(n937), .B(n938), .Y(n515));
sg13g2_inv_4 U916 (.A(last_key_i_116_), .Y(n935));
sg13g2_nand2_2 U917 (.A(n941), .B(n942), .Y(n517));
sg13g2_inv_4 U918 (.A(last_key_i_148_), .Y(n939));
sg13g2_xnor2_1 U919 (.A(last_key_i_84_), .B(n515), .Y(n512));
sg13g2_nor2_2 U920 (.A(n187), .B(round_i_2_), .Y(n131));
sg13g2_nand2_2 U921 (.A(last_key_i_17_), .B(n9), .Y(n36));
sg13g2_xnor2_1 U922 (.A(last_key_i_156_), .B(n125), .Y(n123));
sg13g2_nand2_2 U923 (.A(n78), .B(last_key_i_90_), .Y(n946));
sg13g2_nand2_2 U924 (.A(n946), .B(n947), .Y(n76));
sg13g2_inv_4 U925 (.A(last_key_i_90_), .Y(n944));
sg13g2_nand2_2 U926 (.A(last_key_i_122_), .B(n81), .Y(n950));
sg13g2_nand2_2 U927 (.A(n950), .B(n951), .Y(n78));
sg13g2_inv_4 U928 (.A(last_key_i_122_), .Y(n948));
sg13g2_inv_4 U929 (.A(n81), .Y(n949));
sg13g2_xnor2_1 U930 (.A(last_key_i_58_), .B(n76), .Y(n73));
sg13g2_o21ai_1 U931 (.A1(net25077), .A2(n76), .B1(n77), .Y(n718));
sg13g2_nand2_2 U932 (.A(sbox_data_i_1_), .B(last_key_i_169_), .Y(n954));
sg13g2_nand2_2 U933 (.A(n414), .B(n953), .Y(n955));
sg13g2_nand2_2 U934 (.A(n955), .B(n954), .Y(n273));
sg13g2_inv_4 U935 (.A(last_key_i_169_), .Y(n953));
sg13g2_inv_4 U936 (.A(round_i_2_), .Y(n90));
sg13g2_xnor2_1 U937 (.A(n148), .B(n149), .Y(n145));
sg13g2_inv_4 U938 (.A(net25830), .Y(net25831));
sg13g2_inv_4 U939 (.A(last_key_i_27_), .Y(n956));
sg13g2_inv_4 U940 (.A(n956), .Y(n957));
sg13g2_o21ai_1 U941 (.A1(n234), .A2(net25105), .B1(n235), .Y(n770));
sg13g2_nand4_1 U942 (.A(n111), .B(round_i_3_), .C(n88), .D(round_i_2_), .Y(n109));
sg13g2_nand2_2 U943 (.A(n131), .B(n132), .Y(n70));
sg13g2_inv_4 U944 (.A(round_i_1_), .Y(n111));
sg13g2_nand2_1 U945 (.A(last_key_i_14_), .B(n993), .Y(n990));
sg13g2_nor2_2 U946 (.A(n39), .B(n7), .Y(n38));
sg13g2_a21oi_2 U947 (.A1(last_key_i_28_), .A2(net39266), .B1(n23), .Y(n22));
sg13g2_nand2_1 U948 (.A(last_key_i_13_), .B(n993), .Y(n989));
sg13g2_xnor2_1 U949 (.A(last_key_i_40_), .B(n211), .Y(n226));
sg13g2_xnor2_1 U950 (.A(last_key_i_126_), .B(n161), .Y(n158));
sg13g2_xnor2_1 U951 (.A(last_key_i_62_), .B(n156), .Y(n153));
sg13g2_xnor2_1 U952 (.A(last_key_i_94_), .B(n158), .Y(n156));
sg13g2_inv_4 U953 (.A(last_key_i_10_), .Y(n30));
sg13g2_a21oi_2 U954 (.A1(n5), .A2(last_key_i_29_), .B1(n18), .Y(n17));
sg13g2_nand2_1 U955 (.A(last_key_i_12_), .B(n993), .Y(n986));
sg13g2_xnor2_1 U956 (.A(last_key_i_46_), .B(n193), .Y(n214));
sg13g2_xnor2_1 U957 (.A(n167), .B(n166), .Y(n163));
sg13g2_nand3_1 U958 (.A(n109), .B(n110), .C(n168), .Y(n166));
sg13g2_xnor2_1 U959 (.A(last_key_i_44_), .B(n199), .Y(n218));
sg13g2_nand2_2 U960 (.A(last_key_i_125_), .B(n143), .Y(n960));
sg13g2_nand2_2 U961 (.A(n960), .B(n961), .Y(n140));
sg13g2_inv_4 U962 (.A(last_key_i_125_), .Y(n958));
sg13g2_inv_4 U963 (.A(n143), .Y(n959));
sg13g2_xnor2_1 U964 (.A(n963), .B(n138), .Y(n962));
sg13g2_xnor2_1 U965 (.A(last_key_i_93_), .B(n140), .Y(n138));
sg13g2_nand2_2 U966 (.A(n67), .B(n68), .Y(n966));
sg13g2_nand2_2 U967 (.A(n964), .B(n965), .Y(n967));
sg13g2_nand2_2 U968 (.A(n966), .B(n967), .Y(n64));
sg13g2_inv_4 U969 (.A(n67), .Y(n964));
sg13g2_inv_4 U970 (.A(n68), .Y(n965));
sg13g2_nand2_2 U971 (.A(last_key_i_121_), .B(n62), .Y(n970));
sg13g2_nand2_2 U972 (.A(n970), .B(n971), .Y(n59));
sg13g2_inv_4 U973 (.A(last_key_i_121_), .Y(n968));
sg13g2_inv_4 U974 (.A(n62), .Y(n969));
sg13g2_xnor2_1 U975 (.A(last_key_i_153_), .B(n64), .Y(n62));
sg13g2_xnor2_1 U976 (.A(last_key_i_89_), .B(n59), .Y(n57));
sg13g2_nand2_2 U977 (.A(n974), .B(n99), .Y(n976));
sg13g2_nand2_2 U978 (.A(n975), .B(n976), .Y(n96));
sg13g2_inv_4 U979 (.A(last_key_i_91_), .Y(n974));
sg13g2_xnor2_1 U980 (.A(last_key_i_59_), .B(n96), .Y(n93));
sg13g2_xnor2_1 U981 (.A(last_key_i_155_), .B(n103), .Y(n101));
sg13g2_xnor2_1 U982 (.A(last_key_i_152_), .B(n580), .Y(n577));
sg13g2_xnor2_1 U983 (.A(n582), .B(n583), .Y(n580));
sg13g2_inv_4 U984 (.A(last_key_i_18_), .Y(n977));
sg13g2_xnor2_1 U985 (.A(last_key_i_95_), .B(n177), .Y(n174));
sg13g2_nand2_1 U986 (.A(last_key_i_11_), .B(n993), .Y(n985));
sg13g2_nor2_2 U987 (.A(n90), .B(round_i_3_), .Y(n112));
sg13g2_xnor2_1 U988 (.A(last_key_i_110_), .B(n265), .Y(n233));
sg13g2_xnor2_1 U989 (.A(last_key_i_111_), .B(n267), .Y(n230));
sg13g2_xnor2_1 U990 (.A(col_24_), .B(last_key_i_184_), .Y(n583));
sg13g2_xnor2_1 U991 (.A(last_key_i_76_), .B(n239), .Y(n199));
sg13g2_xnor2_1 U992 (.A(last_key_i_108_), .B(n809), .Y(n239));
sg13g2_xnor2_1 U993 (.A(last_key_i_127_), .B(n179), .Y(n177));
sg13g2_inv_4 U994 (.A(last_key_i_24_), .Y(n978));
sg13g2_inv_4 U995 (.A(last_key_i_29_), .Y(n979));
sg13g2_xnor2_1 U996 (.A(last_key_i_105_), .B(n255), .Y(n248));
sg13g2_xnor2_1 U997 (.A(last_key_i_109_), .B(n263), .Y(n236));
sg13g2_nand2_2 U998 (.A(n982), .B(n983), .Y(n208));
sg13g2_inv_4 U999 (.A(last_key_i_73_), .Y(n980));
sg13g2_inv_4 U1000 (.A(last_key_i_3_), .Y(n29));
sg13g2_xnor2_1 U1001 (.A(last_key_i_107_), .B(n259), .Y(n242));
sg13g2_xnor2_1 U1002 (.A(last_key_i_106_), .B(n257), .Y(n245));
sg13g2_buf_8 U1003 (.A(n52), .X(net25075));
sg13g2_buf_8 U1004 (.A(n52), .X(net25077));
sg13g2_buf_8 U1005 (.A(n52), .X(net25079));
sg13g2_buf_8 U1006 (.A(n52), .X(net25081));
sg13g2_buf_8 U1007 (.A(n52), .X(net25083));
sg13g2_buf_8 U1008 (.A(n52), .X(net25093));
sg13g2_buf_8 U1009 (.A(n52), .X(net25097));
sg13g2_buf_8 U1010 (.A(n52), .X(net25103));
sg13g2_buf_8 U1011 (.A(n52), .X(net25105));
sg13g2_buf_8 U1012 (.A(n52), .X(net25107));
sg13g2_buf_8 U1013 (.A(n52), .X(net25109));
sg13g2_buf_8 U1014 (.A(n52), .X(net25111));
sg13g2_buf_8 U1015 (.A(n52), .X(net25113));
sg13g2_buf_8 U1016 (.A(n52), .X(net25115));
sg13g2_buf_8 U1017 (.A(n52), .X(net25127));
sg13g2_tielo U1018 (.L_LO(sbox_decrypt_o));
sg13g2_nand2_1 U1019 (.A(last_key_i_10_), .B(n993), .Y(n991));
sg13g2_nand2_1 U1020 (.A(n839), .B(n993), .Y(n826));
sg13g2_nand2_1 U1021 (.A(last_key_i_8_), .B(n993), .Y(n987));
sg13g2_dfrbp_1 col_reg_0_ (.CLK(clk), .D(n584), .Q(col_0), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_1_ (.CLK(clk), .D(n585), .Q(col_1), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_2_ (.CLK(clk), .D(n586), .Q(col_2), .RESET_B(reset));
sg13g2_dfrbp_2 col_reg_3_ (.CLK(clk), .D(n587), .Q(col_3), .Q_N(n880), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_4_ (.CLK(clk), .D(n588), .Q(col_4), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_5_ (.CLK(clk), .D(n589), .Q(col_5), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_6_ (.CLK(clk), .D(n590), .Q(col_6), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_7_ (.CLK(clk), .D(n591), .Q(col_7), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_16_ (.CLK(clk), .D(n592), .Q(col_16_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_17_ (.CLK(clk), .D(n593), .Q(col_17_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_18_ (.CLK(clk), .D(n594), .Q(col_18_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_19_ (.CLK(clk), .D(n595), .Q(col_19_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_20_ (.CLK(clk), .D(n596), .Q(col_20_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_21_ (.CLK(clk), .D(n597), .Q(col_21_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_22_ (.CLK(clk), .D(n598), .Q(col_22_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_23_ (.CLK(clk), .D(n599), .Q(col_23_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_24_ (.CLK(clk), .D(n600), .Q(col_24_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_25_ (.CLK(clk), .D(n601), .Q(col_25_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_26_ (.CLK(clk), .D(n602), .Q(col_26_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_27_ (.CLK(clk), .D(n603), .Q(col_27_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_28_ (.CLK(clk), .D(n604), .Q(col_28_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_29_ (.CLK(clk), .D(n605), .Q(col_29_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_30_ (.CLK(clk), .D(n606), .Q(col_30_), .RESET_B(reset));
sg13g2_dfrbp_1 col_reg_31_ (.CLK(clk), .D(n607), .Q(col_31_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_0_ (.CLK(clk), .D(n609), .Q(new_key_o_0_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_1_ (.CLK(clk), .D(n615), .Q(new_key_o_1_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_2_ (.CLK(clk), .D(n621), .Q(new_key_o_2_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_3_ (.CLK(clk), .D(n627), .Q(new_key_o_3_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_4_ (.CLK(clk), .D(n633), .Q(new_key_o_4_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_5_ (.CLK(clk), .D(n639), .Q(new_key_o_5_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_6_ (.CLK(clk), .D(n645), .Q(new_key_o_6_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_7_ (.CLK(clk), .D(n651), .Q(new_key_o_7_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_8_ (.CLK(clk), .D(n775), .Q(new_key_o_8_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_9_ (.CLK(clk), .D(n774), .Q(new_key_o_9_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_10_ (.CLK(clk), .D(n773), .Q(new_key_o_10_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_11_ (.CLK(clk), .D(n772), .Q(new_key_o_11_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_12_ (.CLK(clk), .D(n771), .Q(new_key_o_12_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_13_ (.CLK(clk), .D(n770), .Q(new_key_o_13_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_14_ (.CLK(clk), .D(n769), .Q(new_key_o_14_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_15_ (.CLK(clk), .D(n768), .Q(new_key_o_15_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_16_ (.CLK(clk), .D(n657), .Q(new_key_o_16_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_17_ (.CLK(clk), .D(n663), .Q(new_key_o_17_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_18_ (.CLK(clk), .D(n669), .Q(new_key_o_18_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_19_ (.CLK(clk), .D(n675), .Q(new_key_o_19_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_20_ (.CLK(clk), .D(n681), .Q(new_key_o_20_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_21_ (.CLK(clk), .D(n687), .Q(new_key_o_21_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_22_ (.CLK(clk), .D(n693), .Q(new_key_o_22_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_23_ (.CLK(clk), .D(n699), .Q(new_key_o_23_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_24_ (.CLK(clk), .D(n705), .Q(new_key_o_24_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_25_ (.CLK(clk), .D(n711), .Q(new_key_o_25_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_26_ (.CLK(clk), .D(n717), .Q(new_key_o_26_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_27_ (.CLK(clk), .D(n723), .Q(new_key_o_27_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_28_ (.CLK(clk), .D(n729), .Q(new_key_o_28_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_29_ (.CLK(clk), .D(n735), .Q(new_key_o_29_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_30_ (.CLK(clk), .D(n741), .Q(new_key_o_30_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_31_ (.CLK(clk), .D(n747), .Q(new_key_o_31_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_32_ (.CLK(clk), .D(n608), .Q(new_key_o_32_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_33_ (.CLK(clk), .D(n614), .Q(new_key_o_33_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_34_ (.CLK(clk), .D(n620), .Q(new_key_o_34_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_35_ (.CLK(clk), .D(n626), .Q(new_key_o_35_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_36_ (.CLK(clk), .D(n632), .Q(new_key_o_36_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_37_ (.CLK(clk), .D(n638), .Q(new_key_o_37_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_38_ (.CLK(clk), .D(n644), .Q(new_key_o_38_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_39_ (.CLK(clk), .D(n650), .Q(new_key_o_39_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_40_ (.CLK(clk), .D(n767), .Q(new_key_o_40_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_41_ (.CLK(clk), .D(n766), .Q(new_key_o_41_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_42_ (.CLK(clk), .D(n765), .Q(new_key_o_42_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_43_ (.CLK(clk), .D(n764), .Q(new_key_o_43_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_44_ (.CLK(clk), .D(n763), .Q(new_key_o_44_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_45_ (.CLK(clk), .D(n762), .Q(new_key_o_45_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_46_ (.CLK(clk), .D(n761), .Q(new_key_o_46_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_47_ (.CLK(clk), .D(n760), .Q(new_key_o_47_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_48_ (.CLK(clk), .D(n656), .Q(new_key_o_48_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_49_ (.CLK(clk), .D(n662), .Q(new_key_o_49_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_50_ (.CLK(clk), .D(n668), .Q(new_key_o_50_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_51_ (.CLK(clk), .D(n674), .Q(new_key_o_51_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_52_ (.CLK(clk), .D(n680), .Q(new_key_o_52_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_53_ (.CLK(clk), .D(n686), .Q(new_key_o_53_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_54_ (.CLK(clk), .D(n692), .Q(new_key_o_54_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_55_ (.CLK(clk), .D(n698), .Q(new_key_o_55_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_56_ (.CLK(clk), .D(n704), .Q(new_key_o_56_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_57_ (.CLK(clk), .D(n710), .Q(new_key_o_57_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_58_ (.CLK(clk), .D(n716), .Q(new_key_o_58_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_59_ (.CLK(clk), .D(n722), .Q(new_key_o_59_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_60_ (.CLK(clk), .D(n728), .Q(new_key_o_60_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_61_ (.CLK(clk), .D(n734), .Q(new_key_o_61_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_62_ (.CLK(clk), .D(n740), .Q(new_key_o_62_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_63_ (.CLK(clk), .D(n746), .Q(new_key_o_63_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_64_ (.CLK(clk), .D(n610), .Q(new_key_o_64_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_65_ (.CLK(clk), .D(n616), .Q(new_key_o_65_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_66_ (.CLK(clk), .D(n622), .Q(new_key_o_66_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_67_ (.CLK(clk), .D(n628), .Q(new_key_o_67_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_68_ (.CLK(clk), .D(n634), .Q(new_key_o_68_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_69_ (.CLK(clk), .D(n640), .Q(new_key_o_69_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_70_ (.CLK(clk), .D(n646), .Q(new_key_o_70_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_71_ (.CLK(clk), .D(n652), .Q(new_key_o_71_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_72_ (.CLK(clk), .D(n759), .Q(new_key_o_72_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_73_ (.CLK(clk), .D(n758), .Q(new_key_o_73_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_74_ (.CLK(clk), .D(n757), .Q(new_key_o_74_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_75_ (.CLK(clk), .D(n756), .Q(new_key_o_75_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_76_ (.CLK(clk), .D(n755), .Q(new_key_o_76_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_77_ (.CLK(clk), .D(n754), .Q(new_key_o_77_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_78_ (.CLK(clk), .D(n753), .Q(new_key_o_78_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_79_ (.CLK(clk), .D(n752), .Q(new_key_o_79_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_80_ (.CLK(clk), .D(n658), .Q(new_key_o_80_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_81_ (.CLK(clk), .D(n664), .Q(new_key_o_81_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_82_ (.CLK(clk), .D(n670), .Q(new_key_o_82_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_83_ (.CLK(clk), .D(n676), .Q(new_key_o_83_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_84_ (.CLK(clk), .D(n682), .Q(new_key_o_84_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_85_ (.CLK(clk), .D(n688), .Q(new_key_o_85_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_86_ (.CLK(clk), .D(n694), .Q(new_key_o_86_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_87_ (.CLK(clk), .D(n700), .Q(new_key_o_87_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_88_ (.CLK(clk), .D(n706), .Q(new_key_o_88_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_89_ (.CLK(clk), .D(n712), .Q(new_key_o_89_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_90_ (.CLK(clk), .D(n718), .Q(new_key_o_90_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_91_ (.CLK(clk), .D(n724), .Q(new_key_o_91_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_92_ (.CLK(clk), .D(n730), .Q(new_key_o_92_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_93_ (.CLK(clk), .D(n736), .Q(new_key_o_93_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_94_ (.CLK(clk), .D(n742), .Q(new_key_o_94_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_95_ (.CLK(clk), .D(n748), .Q(new_key_o_95_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_96_ (.CLK(clk), .D(n611), .Q(new_key_o_96_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_97_ (.CLK(clk), .D(n617), .Q(new_key_o_97_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_98_ (.CLK(clk), .D(n623), .Q(new_key_o_98_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_99_ (.CLK(clk), .D(n629), .Q(new_key_o_99_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_100_ (.CLK(clk), .D(n635), .Q(new_key_o_100_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_101_ (.CLK(clk), .D(n641), .Q(new_key_o_101_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_102_ (.CLK(clk), .D(n647), .Q(new_key_o_102_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_103_ (.CLK(clk), .D(n653), .Q(new_key_o_103_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_104_ (.CLK(clk), .D(n776), .Q(new_key_o_104_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_105_ (.CLK(clk), .D(n777), .Q(new_key_o_105_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_106_ (.CLK(clk), .D(n778), .Q(new_key_o_106_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_107_ (.CLK(clk), .D(n779), .Q(new_key_o_107_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_108_ (.CLK(clk), .D(n780), .Q(new_key_o_108_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_109_ (.CLK(clk), .D(n781), .Q(new_key_o_109_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_110_ (.CLK(clk), .D(n782), .Q(new_key_o_110_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_111_ (.CLK(clk), .D(n783), .Q(new_key_o_111_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_112_ (.CLK(clk), .D(n659), .Q(new_key_o_112_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_113_ (.CLK(clk), .D(n665), .Q(new_key_o_113_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_114_ (.CLK(clk), .D(n671), .Q(new_key_o_114_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_115_ (.CLK(clk), .D(n677), .Q(new_key_o_115_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_116_ (.CLK(clk), .D(n683), .Q(new_key_o_116_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_117_ (.CLK(clk), .D(n689), .Q(new_key_o_117_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_118_ (.CLK(clk), .D(n695), .Q(new_key_o_118_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_119_ (.CLK(clk), .D(n701), .Q(new_key_o_119_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_120_ (.CLK(clk), .D(n707), .Q(new_key_o_120_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_121_ (.CLK(clk), .D(n713), .Q(new_key_o_121_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_122_ (.CLK(clk), .D(n719), .Q(new_key_o_122_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_123_ (.CLK(clk), .D(n725), .Q(new_key_o_123_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_124_ (.CLK(clk), .D(n731), .Q(new_key_o_124_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_125_ (.CLK(clk), .D(n737), .Q(new_key_o_125_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_126_ (.CLK(clk), .D(n743), .Q(new_key_o_126_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_127_ (.CLK(clk), .D(n749), .Q(new_key_o_127_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_128_ (.CLK(clk), .D(n612), .Q(new_key_o_128_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_129_ (.CLK(clk), .D(n618), .Q(new_key_o_129_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_130_ (.CLK(clk), .D(n624), .Q(new_key_o_130_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_131_ (.CLK(clk), .D(n630), .Q(new_key_o_131_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_132_ (.CLK(clk), .D(n636), .Q(new_key_o_132_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_133_ (.CLK(clk), .D(n642), .Q(new_key_o_133_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_134_ (.CLK(clk), .D(n648), .Q(new_key_o_134_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_135_ (.CLK(clk), .D(n654), .Q(new_key_o_135_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_136_ (.CLK(clk), .D(n784), .Q(new_key_o_136_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_137_ (.CLK(clk), .D(n785), .Q(new_key_o_137_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_138_ (.CLK(clk), .D(n786), .Q(new_key_o_138_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_139_ (.CLK(clk), .D(n787), .Q(new_key_o_139_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_140_ (.CLK(clk), .D(n788), .Q(new_key_o_140_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_141_ (.CLK(clk), .D(n789), .Q(new_key_o_141_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_142_ (.CLK(clk), .D(n790), .Q(new_key_o_142_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_143_ (.CLK(clk), .D(n791), .Q(new_key_o_143_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_144_ (.CLK(clk), .D(n660), .Q(new_key_o_144_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_145_ (.CLK(clk), .D(n666), .Q(new_key_o_145_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_146_ (.CLK(clk), .D(n672), .Q(new_key_o_146_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_147_ (.CLK(clk), .D(n678), .Q(new_key_o_147_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_148_ (.CLK(clk), .D(n684), .Q(new_key_o_148_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_149_ (.CLK(clk), .D(n690), .Q(new_key_o_149_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_150_ (.CLK(clk), .D(n696), .Q(new_key_o_150_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_151_ (.CLK(clk), .D(n702), .Q(new_key_o_151_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_152_ (.CLK(clk), .D(n708), .Q(new_key_o_152_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_153_ (.CLK(clk), .D(n714), .Q(new_key_o_153_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_154_ (.CLK(clk), .D(n720), .Q(new_key_o_154_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_155_ (.CLK(clk), .D(n726), .Q(new_key_o_155_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_156_ (.CLK(clk), .D(n732), .Q(new_key_o_156_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_157_ (.CLK(clk), .D(n738), .Q(new_key_o_157_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_158_ (.CLK(clk), .D(n744), .Q(new_key_o_158_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_159_ (.CLK(clk), .D(n750), .Q(new_key_o_159_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_160_ (.CLK(clk), .D(n613), .Q(new_key_o_160_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_161_ (.CLK(clk), .D(n619), .Q(new_key_o_161_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_162_ (.CLK(clk), .D(n625), .Q(new_key_o_162_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_163_ (.CLK(clk), .D(n631), .Q(new_key_o_163_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_164_ (.CLK(clk), .D(n637), .Q(new_key_o_164_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_165_ (.CLK(clk), .D(n643), .Q(new_key_o_165_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_166_ (.CLK(clk), .D(n649), .Q(new_key_o_166_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_167_ (.CLK(clk), .D(n655), .Q(new_key_o_167_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_168_ (.CLK(clk), .D(n792), .Q(new_key_o_168_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_169_ (.CLK(clk), .D(n793), .Q(new_key_o_169_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_170_ (.CLK(clk), .D(n794), .Q(new_key_o_170_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_171_ (.CLK(clk), .D(n795), .Q(new_key_o_171_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_172_ (.CLK(clk), .D(n796), .Q(new_key_o_172_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_173_ (.CLK(clk), .D(n797), .Q(new_key_o_173_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_174_ (.CLK(clk), .D(n798), .Q(new_key_o_174_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_175_ (.CLK(clk), .D(n799), .Q(new_key_o_175_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_176_ (.CLK(clk), .D(n661), .Q(new_key_o_176_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_177_ (.CLK(clk), .D(n667), .Q(new_key_o_177_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_178_ (.CLK(clk), .D(n673), .Q(new_key_o_178_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_179_ (.CLK(clk), .D(n679), .Q(new_key_o_179_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_180_ (.CLK(clk), .D(n685), .Q(new_key_o_180_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_181_ (.CLK(clk), .D(n691), .Q(new_key_o_181_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_182_ (.CLK(clk), .D(n697), .Q(new_key_o_182_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_183_ (.CLK(clk), .D(n703), .Q(new_key_o_183_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_184_ (.CLK(clk), .D(n709), .Q(new_key_o_184_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_185_ (.CLK(clk), .D(n715), .Q(new_key_o_185_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_186_ (.CLK(clk), .D(n721), .Q(new_key_o_186_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_187_ (.CLK(clk), .D(n727), .Q(new_key_o_187_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_188_ (.CLK(clk), .D(n733), .Q(new_key_o_188_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_189_ (.CLK(clk), .D(n739), .Q(new_key_o_189_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_190_ (.CLK(clk), .D(n745), .Q(new_key_o_190_), .RESET_B(reset));
sg13g2_dfrbp_1 key_reg_reg_191_ (.CLK(clk), .D(n751), .Q(new_key_o_191_), .RESET_B(reset));
sg13g2_dfrbp_1 ready_o_reg (.CLK(clk), .D(next_ready_o), .Q(ready_o), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_0_ (.CLK(clk), .D(n801), .Q(state_0_), .Q_N(n49), .RESET_B(reset));
sg13g2_dfrbp_1 state_reg_1_ (.CLK(clk), .D(n800), .Q(state_1_), .Q_N(n50), .RESET_B(reset));
sg13g2_dfrbp_2 state_reg_2_ (.CLK(clk), .D(n855), .Q(state_2_), .Q_N(n318), .RESET_B(reset));
endmodule

