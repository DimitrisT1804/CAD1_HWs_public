// Generated netlist by CADI API on Date: 2025-10-23 15:02:51 //

module PID_1 (\i_wb_adr[0], \i_wb_adr[1], \i_wb_adr[2], \i_wb_adr[3], \i_wb_adr[4], \i_wb_adr[5], \i_wb_adr[6], \i_wb_adr[7], \i_wb_adr[8], \i_wb_adr[9], \i_wb_adr[10], \i_wb_adr[11], \i_wb_adr[12], \i_wb_adr[13], \i_wb_adr[14], \i_wb_adr[15], \i_wb_data[0], \i_wb_data[1], \i_wb_data[2], \i_wb_data[3], \i_wb_data[4], \i_wb_data[5], \i_wb_data[6], \i_wb_data[7], \i_wb_data[8], \i_wb_data[9], \i_wb_data[10], \i_wb_data[11], \i_wb_data[12], \i_wb_data[13], \i_wb_data[14], \i_wb_data[15], \i_wb_data[16], \i_wb_data[17], \i_wb_data[18], \i_wb_data[19], \i_wb_data[20], \i_wb_data[21], \i_wb_data[22], \i_wb_data[23], \i_wb_data[24], \i_wb_data[25], \i_wb_data[26], \i_wb_data[27], \i_wb_data[28], \i_wb_data[29], \i_wb_data[30], \i_wb_data[31], \o_un[0], \o_un[1], \o_un[2], \o_un[3], \o_un[4], \o_un[5], \o_un[6], \o_un[7], \o_un[8], \o_un[9], \o_un[10], \o_un[11], \o_un[12], \o_un[13], \o_un[14], \o_un[15], \o_un[16], \o_un[17], \o_un[18], \o_un[19], \o_un[20], \o_un[21], \o_un[22], \o_un[23], \o_un[24], \o_un[25], \o_un[26], \o_un[27], \o_un[28], \o_un[29], \o_un[30], \o_un[31], \o_wb_data[0], \o_wb_data[1], \o_wb_data[2], \o_wb_data[3], \o_wb_data[4], \o_wb_data[5], \o_wb_data[6], \o_wb_data[7], \o_wb_data[8], \o_wb_data[9], \o_wb_data[10], \o_wb_data[11], \o_wb_data[12], \o_wb_data[13], \o_wb_data[14], \o_wb_data[15], \o_wb_data[16], \o_wb_data[17], \o_wb_data[18], \o_wb_data[19], \o_wb_data[20], \o_wb_data[21], \o_wb_data[22], \o_wb_data[23], \o_wb_data[24], \o_wb_data[25], \o_wb_data[26], \o_wb_data[27], \o_wb_data[28], \o_wb_data[29], \o_wb_data[30], \o_wb_data[31], i_clk, i_rst, i_wb_cyc, i_wb_stb, i_wb_we, o_valid, o_wb_ack);
input \i_wb_adr[0], \i_wb_adr[1], \i_wb_adr[2], \i_wb_adr[3], \i_wb_adr[4], \i_wb_adr[5], \i_wb_adr[6], \i_wb_adr[7], \i_wb_adr[8], \i_wb_adr[9], \i_wb_adr[10], \i_wb_adr[11], \i_wb_adr[12], \i_wb_adr[13], \i_wb_adr[14], \i_wb_adr[15], \i_wb_data[0], \i_wb_data[1], \i_wb_data[2], \i_wb_data[3], \i_wb_data[4], \i_wb_data[5], \i_wb_data[6], \i_wb_data[7], \i_wb_data[8], \i_wb_data[9], \i_wb_data[10], \i_wb_data[11], \i_wb_data[12], \i_wb_data[13], \i_wb_data[14], \i_wb_data[15], \i_wb_data[16], \i_wb_data[17], \i_wb_data[18], \i_wb_data[19], \i_wb_data[20], \i_wb_data[21], \i_wb_data[22], \i_wb_data[23], \i_wb_data[24], \i_wb_data[25], \i_wb_data[26], \i_wb_data[27], \i_wb_data[28], \i_wb_data[29], \i_wb_data[30], \i_wb_data[31], i_clk, i_rst, i_wb_cyc, i_wb_stb, i_wb_we;
output \o_un[0], \o_un[1], \o_un[2], \o_un[3], \o_un[4], \o_un[5], \o_un[6], \o_un[7], \o_un[8], \o_un[9], \o_un[10], \o_un[11], \o_un[12], \o_un[13], \o_un[14], \o_un[15], \o_un[16], \o_un[17], \o_un[18], \o_un[19], \o_un[20], \o_un[21], \o_un[22], \o_un[23], \o_un[24], \o_un[25], \o_un[26], \o_un[27], \o_un[28], \o_un[29], \o_un[30], \o_un[31], \o_wb_data[0], \o_wb_data[1], \o_wb_data[2], \o_wb_data[3], \o_wb_data[4], \o_wb_data[5], \o_wb_data[6], \o_wb_data[7], \o_wb_data[8], \o_wb_data[9], \o_wb_data[10], \o_wb_data[11], \o_wb_data[12], \o_wb_data[13], \o_wb_data[14], \o_wb_data[15], \o_wb_data[16], \o_wb_data[17], \o_wb_data[18], \o_wb_data[19], \o_wb_data[20], \o_wb_data[21], \o_wb_data[22], \o_wb_data[23], \o_wb_data[24], \o_wb_data[25], \o_wb_data[26], \o_wb_data[27], \o_wb_data[28], \o_wb_data[29], \o_wb_data[30], \o_wb_data[31], o_valid, o_wb_ack;

sg13g2_dfrbp_1 \a_reg[0] (.CLK(i_clk), .D(n876), .Q(a_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[1] (.CLK(i_clk), .D(n875), .Q(a_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[2] (.CLK(i_clk), .D(n874), .Q(a_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[3] (.CLK(i_clk), .D(n873), .Q(a_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[4] (.CLK(i_clk), .D(n872), .Q(a_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[5] (.CLK(i_clk), .D(n871), .Q(a_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[6] (.CLK(i_clk), .D(n870), .Q(a_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[7] (.CLK(i_clk), .D(n869), .Q(a_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[8] (.CLK(i_clk), .D(n868), .Q(a_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[9] (.CLK(i_clk), .D(n867), .Q(a_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[10] (.CLK(i_clk), .D(n866), .Q(a_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[11] (.CLK(i_clk), .D(n865), .Q(a_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[12] (.CLK(i_clk), .D(n864), .Q(a_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[13] (.CLK(i_clk), .D(n863), .Q(a_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[14] (.CLK(i_clk), .D(n862), .Q(a_14), .RESET_B(n1340));
sg13g2_dfrbp_2 \a_reg[15] (.CLK(i_clk), .D(n861), .Q(a_15), .Q_N(N551), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[16] (.CLK(i_clk), .D(n857), .Q(a_16), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[17] (.CLK(i_clk), .D(n856), .Q(a_17), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[18] (.CLK(i_clk), .D(n855), .Q(a_18), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[19] (.CLK(i_clk), .D(n854), .Q(a_19), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[20] (.CLK(i_clk), .D(n853), .Q(a_20), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[21] (.CLK(i_clk), .D(n852), .Q(a_21), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[22] (.CLK(i_clk), .D(n851), .Q(a_22), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[23] (.CLK(i_clk), .D(n850), .Q(a_23), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[24] (.CLK(i_clk), .D(n849), .Q(a_24), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[25] (.CLK(i_clk), .D(n848), .Q(a_25), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[26] (.CLK(i_clk), .D(n847), .Q(a_26), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[27] (.CLK(i_clk), .D(n846), .Q(a_27), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[28] (.CLK(i_clk), .D(n845), .Q(a_28), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[29] (.CLK(i_clk), .D(n844), .Q(a_29), .RESET_B(n1340));
sg13g2_dfrbp_1 \a_reg[30] (.CLK(i_clk), .D(n843), .Q(a_30), .RESET_B(n1340));
sg13g2_dfrbp_2 \a_reg[31] (.CLK(i_clk), .D(n842), .Q(a_31), .Q_N(N558), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][0] (.CLK(i_clk), .D(n956), .Q(\err[0][0]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][1] (.CLK(i_clk), .D(n955), .Q(\err[0][1]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][2] (.CLK(i_clk), .D(n954), .Q(\err[0][2]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][3] (.CLK(i_clk), .D(n953), .Q(\err[0][3]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][4] (.CLK(i_clk), .D(n952), .Q(\err[0][4]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][5] (.CLK(i_clk), .D(n951), .Q(\err[0][5]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][6] (.CLK(i_clk), .D(n950), .Q(\err[0][6]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][7] (.CLK(i_clk), .D(n949), .Q(\err[0][7]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][8] (.CLK(i_clk), .D(n948), .Q(\err[0][8]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][9] (.CLK(i_clk), .D(n947), .Q(\err[0][9]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][10] (.CLK(i_clk), .D(n946), .Q(\err[0][10]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][11] (.CLK(i_clk), .D(n945), .Q(\err[0][11]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][12] (.CLK(i_clk), .D(n944), .Q(\err[0][12]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][13] (.CLK(i_clk), .D(n943), .Q(\err[0][13]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][14] (.CLK(i_clk), .D(n942), .Q(\err[0][14]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[0][15] (.CLK(i_clk), .D(n941), .Q(\err[0][15]), .Q_N(n422), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][0] (.CLK(i_clk), .D(n34), .Q(\err[1][0]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][1] (.CLK(i_clk), .D(n33), .Q(\err[1][1]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][2] (.CLK(i_clk), .D(n32), .Q(\err[1][2]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][3] (.CLK(i_clk), .D(n31), .Q(\err[1][3]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][4] (.CLK(i_clk), .D(n30), .Q(\err[1][4]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][5] (.CLK(i_clk), .D(n29), .Q(\err[1][5]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][6] (.CLK(i_clk), .D(n28), .Q(\err[1][6]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][7] (.CLK(i_clk), .D(n27), .Q(\err[1][7]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][8] (.CLK(i_clk), .D(n26), .Q(\err[1][8]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][9] (.CLK(i_clk), .D(n25), .Q(\err[1][9]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][10] (.CLK(i_clk), .D(n24), .Q(\err[1][10]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][11] (.CLK(i_clk), .D(n23), .Q(\err[1][11]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][12] (.CLK(i_clk), .D(n22), .Q(\err[1][12]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][13] (.CLK(i_clk), .D(n21), .Q(\err[1][13]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][14] (.CLK(i_clk), .D(n20), .Q(\err[1][14]), .RESET_B(n1340));
sg13g2_dfrbp_1 \err_reg[1][15] (.CLK(i_clk), .D(n19), .Q(\err[1][15]), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[0] (.CLK(i_clk), .D(n1087), .Q(kd_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[1] (.CLK(i_clk), .D(n1086), .Q(kd_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[2] (.CLK(i_clk), .D(n1085), .Q(kd_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[3] (.CLK(i_clk), .D(n1084), .Q(kd_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[4] (.CLK(i_clk), .D(n1083), .Q(kd_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[5] (.CLK(i_clk), .D(n1082), .Q(kd_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[6] (.CLK(i_clk), .D(n1081), .Q(kd_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[7] (.CLK(i_clk), .D(n1080), .Q(kd_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[8] (.CLK(i_clk), .D(n1079), .Q(kd_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[9] (.CLK(i_clk), .D(n1078), .Q(kd_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[10] (.CLK(i_clk), .D(n1077), .Q(kd_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[11] (.CLK(i_clk), .D(n1076), .Q(kd_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[12] (.CLK(i_clk), .D(n1075), .Q(kd_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[13] (.CLK(i_clk), .D(n1074), .Q(kd_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[14] (.CLK(i_clk), .D(n1073), .Q(kd_14), .RESET_B(n1340));
sg13g2_dfrbp_1 \kd_reg[15] (.CLK(i_clk), .D(n1072), .Q(kd_15), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[0] (.CLK(i_clk), .D(n1103), .Q(ki_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[1] (.CLK(i_clk), .D(n1102), .Q(ki_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[2] (.CLK(i_clk), .D(n1101), .Q(ki_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[3] (.CLK(i_clk), .D(n1100), .Q(ki_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[4] (.CLK(i_clk), .D(n1099), .Q(ki_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[5] (.CLK(i_clk), .D(n1098), .Q(ki_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[6] (.CLK(i_clk), .D(n1097), .Q(ki_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[7] (.CLK(i_clk), .D(n1096), .Q(ki_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[8] (.CLK(i_clk), .D(n1095), .Q(ki_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[9] (.CLK(i_clk), .D(n1094), .Q(ki_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[10] (.CLK(i_clk), .D(n1093), .Q(ki_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[11] (.CLK(i_clk), .D(n1092), .Q(ki_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[12] (.CLK(i_clk), .D(n1091), .Q(ki_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[13] (.CLK(i_clk), .D(n1090), .Q(ki_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[14] (.CLK(i_clk), .D(n1089), .Q(ki_14), .RESET_B(n1340));
sg13g2_dfrbp_1 \ki_reg[15] (.CLK(i_clk), .D(n1088), .Q(ki_15), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[0] (.CLK(i_clk), .D(n1039), .Q(kp_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[1] (.CLK(i_clk), .D(n1038), .Q(kp_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[2] (.CLK(i_clk), .D(n1037), .Q(kp_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[3] (.CLK(i_clk), .D(n1036), .Q(kp_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[4] (.CLK(i_clk), .D(n1035), .Q(kp_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[5] (.CLK(i_clk), .D(n1034), .Q(kp_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[6] (.CLK(i_clk), .D(n1033), .Q(kp_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[7] (.CLK(i_clk), .D(n1032), .Q(kp_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[8] (.CLK(i_clk), .D(n1031), .Q(kp_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[9] (.CLK(i_clk), .D(n1030), .Q(kp_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[10] (.CLK(i_clk), .D(n1029), .Q(kp_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[11] (.CLK(i_clk), .D(n1028), .Q(kp_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[12] (.CLK(i_clk), .D(n1027), .Q(kp_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[13] (.CLK(i_clk), .D(n1026), .Q(kp_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[14] (.CLK(i_clk), .D(n1025), .Q(kp_14), .RESET_B(n1340));
sg13g2_dfrbp_1 \kp_reg[15] (.CLK(i_clk), .D(n1024), .Q(kp_15), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[0] (.CLK(i_clk), .D(n972), .Q(kpd_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[1] (.CLK(i_clk), .D(n971), .Q(kpd_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[2] (.CLK(i_clk), .D(n970), .Q(kpd_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[3] (.CLK(i_clk), .D(n969), .Q(kpd_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[4] (.CLK(i_clk), .D(n968), .Q(kpd_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[5] (.CLK(i_clk), .D(n967), .Q(kpd_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[6] (.CLK(i_clk), .D(n966), .Q(kpd_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[7] (.CLK(i_clk), .D(n965), .Q(kpd_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[8] (.CLK(i_clk), .D(n964), .Q(kpd_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[9] (.CLK(i_clk), .D(n963), .Q(kpd_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[10] (.CLK(i_clk), .D(n962), .Q(kpd_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[11] (.CLK(i_clk), .D(n961), .Q(kpd_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[12] (.CLK(i_clk), .D(n960), .Q(kpd_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[13] (.CLK(i_clk), .D(n959), .Q(kpd_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[14] (.CLK(i_clk), .D(n958), .Q(kpd_14), .RESET_B(n1340));
sg13g2_dfrbp_1 \kpd_reg[15] (.CLK(i_clk), .D(n957), .Q(kpd_15), .RESET_B(n1340));
sg13g2_dfrbp_1 \md_index_reg[0] (.CLK(i_clk), .D(n1005), .Q(md_index_0), .Q_N(n1248), .RESET_B(n1340));
sg13g2_dfrbp_1 \md_index_reg[1] (.CLK(i_clk), .D(n1006), .Q(md_index_1), .Q_N(n1251), .RESET_B(n1340));
sg13g2_dfrbp_2 \mr_index_reg[0] (.CLK(i_clk), .D(n1007), .Q(mr_index_0), .Q_N(N474), .RESET_B(n1340));
sg13g2_dfrbp_1 \mr_index_reg[1] (.CLK(i_clk), .D(n1008), .Q(mr_index_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \of_reg[0] (.CLK(i_clk), .D(n858), .Q(of_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \of_reg[1] (.CLK(i_clk), .D(n860), .Q(of_1), .Q_N(n379), .RESET_B(n1340));
sg13g2_dfrbp_1 \of_reg[2] (.CLK(i_clk), .D(n859), .Q(of_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \of_reg[3] (.CLK(i_clk), .D(n840), .Q(of_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \of_reg[4] (.CLK(i_clk), .D(n841), .Q(of_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[0] (.CLK(i_clk), .D(n1004), .Q(p_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[1] (.CLK(i_clk), .D(n1003), .Q(p_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[2] (.CLK(i_clk), .D(n1002), .Q(p_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[3] (.CLK(i_clk), .D(n1001), .Q(p_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[4] (.CLK(i_clk), .D(n1000), .Q(p_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[5] (.CLK(i_clk), .D(n999), .Q(p_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[6] (.CLK(i_clk), .D(n998), .Q(p_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[7] (.CLK(i_clk), .D(n997), .Q(p_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[8] (.CLK(i_clk), .D(n996), .Q(p_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[9] (.CLK(i_clk), .D(n995), .Q(p_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[10] (.CLK(i_clk), .D(n994), .Q(p_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[11] (.CLK(i_clk), .D(n993), .Q(p_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[12] (.CLK(i_clk), .D(n992), .Q(p_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[13] (.CLK(i_clk), .D(n991), .Q(p_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[14] (.CLK(i_clk), .D(n990), .Q(p_14), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[15] (.CLK(i_clk), .D(n989), .Q(p_15), .Q_N(N550), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[16] (.CLK(i_clk), .D(n988), .Q(p_16), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[17] (.CLK(i_clk), .D(n987), .Q(p_17), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[18] (.CLK(i_clk), .D(n986), .Q(p_18), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[19] (.CLK(i_clk), .D(n1300), .Q(p_19), .Q_N(n1299), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[20] (.CLK(i_clk), .D(n1305), .Q(p_20), .Q_N(n1304), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[21] (.CLK(i_clk), .D(n983), .Q(p_21), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[22] (.CLK(i_clk), .D(n1327), .Q(p_22), .Q_N(n1328), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[23] (.CLK(i_clk), .D(n981), .Q(p_23), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[24] (.CLK(i_clk), .D(n980), .Q(p_24), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[25] (.CLK(i_clk), .D(n979), .Q(p_25), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[26] (.CLK(i_clk), .D(n978), .Q(p_26), .RESET_B(n1340));
sg13g2_dfrbp_1 \p_reg[27] (.CLK(i_clk), .D(n977), .Q(p_27), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[28] (.CLK(i_clk), .D(n1311), .Q(p_28), .Q_N(n1312), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[29] (.CLK(i_clk), .D(n1325), .Q(p_29), .Q_N(n1326), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[30] (.CLK(i_clk), .D(net9912), .Q(p_30), .Q_N(net9913), .RESET_B(n1340));
sg13g2_dfrbp_2 \p_reg[31] (.CLK(i_clk), .D(n1309), .Q(p_31), .Q_N(N557), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[0] (.CLK(i_clk), .D(n1055), .Q(pv_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[1] (.CLK(i_clk), .D(n1054), .Q(pv_1), .Q_N(n424), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[2] (.CLK(i_clk), .D(n1053), .Q(pv_2), .Q_N(n435), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[3] (.CLK(i_clk), .D(n1052), .Q(pv_3), .Q_N(n442), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[4] (.CLK(i_clk), .D(n1051), .Q(pv_4), .Q_N(n436), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[5] (.CLK(i_clk), .D(n1050), .Q(pv_5), .Q_N(n437), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[6] (.CLK(i_clk), .D(n1049), .Q(pv_6), .Q_N(n438), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[7] (.CLK(i_clk), .D(n1048), .Q(pv_7), .Q_N(n439), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[8] (.CLK(i_clk), .D(n1047), .Q(pv_8), .Q_N(n428), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[9] (.CLK(i_clk), .D(n1046), .Q(pv_9), .Q_N(n434), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[10] (.CLK(i_clk), .D(n1045), .Q(pv_10), .Q_N(n425), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[11] (.CLK(i_clk), .D(n1044), .Q(pv_11), .Q_N(n433), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[12] (.CLK(i_clk), .D(n1043), .Q(pv_12), .Q_N(n441), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[13] (.CLK(i_clk), .D(n1042), .Q(pv_13), .Q_N(n440), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[14] (.CLK(i_clk), .D(n1041), .Q(pv_14), .Q_N(n427), .RESET_B(n1340));
sg13g2_dfrbp_1 \pv_reg[15] (.CLK(i_clk), .D(n1040), .Q(pv_15), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[0] (.CLK(i_clk), .D(n908), .Q(sigma_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[1] (.CLK(i_clk), .D(n907), .Q(sigma_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[2] (.CLK(i_clk), .D(n906), .Q(sigma_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[3] (.CLK(i_clk), .D(n905), .Q(sigma_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[4] (.CLK(i_clk), .D(n904), .Q(sigma_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[5] (.CLK(i_clk), .D(n903), .Q(sigma_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[6] (.CLK(i_clk), .D(n902), .Q(sigma_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[7] (.CLK(i_clk), .D(n901), .Q(sigma_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[8] (.CLK(i_clk), .D(n900), .Q(sigma_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[9] (.CLK(i_clk), .D(n899), .Q(sigma_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[10] (.CLK(i_clk), .D(n898), .Q(sigma_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[11] (.CLK(i_clk), .D(n897), .Q(sigma_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[12] (.CLK(i_clk), .D(n896), .Q(sigma_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[13] (.CLK(i_clk), .D(n895), .Q(sigma_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[14] (.CLK(i_clk), .D(n894), .Q(sigma_14), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[15] (.CLK(i_clk), .D(n893), .Q(sigma_15), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[16] (.CLK(i_clk), .D(n892), .Q(sigma_16), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[17] (.CLK(i_clk), .D(n891), .Q(sigma_17), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[18] (.CLK(i_clk), .D(n890), .Q(sigma_18), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[19] (.CLK(i_clk), .D(n889), .Q(sigma_19), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[20] (.CLK(i_clk), .D(n888), .Q(sigma_20), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[21] (.CLK(i_clk), .D(n887), .Q(sigma_21), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[22] (.CLK(i_clk), .D(n886), .Q(sigma_22), .Q_N(n1306), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[23] (.CLK(i_clk), .D(n885), .Q(sigma_23), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[24] (.CLK(i_clk), .D(n884), .Q(sigma_24), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[25] (.CLK(i_clk), .D(n883), .Q(sigma_25), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[26] (.CLK(i_clk), .D(n882), .Q(sigma_26), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[27] (.CLK(i_clk), .D(n881), .Q(sigma_27), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[28] (.CLK(i_clk), .D(n880), .Q(sigma_28), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[29] (.CLK(i_clk), .D(n879), .Q(sigma_29), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[30] (.CLK(i_clk), .D(n878), .Q(sigma_30), .RESET_B(n1340));
sg13g2_dfrbp_1 \sigma_reg[31] (.CLK(i_clk), .D(n877), .Q(sigma_31), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[0] (.CLK(i_clk), .D(n1071), .Q(sp_0), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[1] (.CLK(i_clk), .D(n1070), .Q(sp_1), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[2] (.CLK(i_clk), .D(n1069), .Q(sp_2), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[3] (.CLK(i_clk), .D(n1068), .Q(sp_3), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[4] (.CLK(i_clk), .D(n1067), .Q(sp_4), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[5] (.CLK(i_clk), .D(n1066), .Q(sp_5), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[6] (.CLK(i_clk), .D(n1065), .Q(sp_6), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[7] (.CLK(i_clk), .D(n1064), .Q(sp_7), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[8] (.CLK(i_clk), .D(n1063), .Q(sp_8), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[9] (.CLK(i_clk), .D(n1062), .Q(sp_9), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[10] (.CLK(i_clk), .D(n1061), .Q(sp_10), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[11] (.CLK(i_clk), .D(n1060), .Q(sp_11), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[12] (.CLK(i_clk), .D(n1059), .Q(sp_12), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[13] (.CLK(i_clk), .D(n1058), .Q(sp_13), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[14] (.CLK(i_clk), .D(n1057), .Q(sp_14), .RESET_B(n1340));
sg13g2_dfrbp_1 \sp_reg[15] (.CLK(i_clk), .D(n1056), .Q(sp_15), .RESET_B(n1340));
sg13g2_sdfbbp_1 \state_1_reg[0] (.CLK(i_clk), .D(n652), .Q(state_1_0), .RESET_B(n1340), .SCD(n651), .SCE(n651), .SET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[1] (.CLK(i_clk), .D(n1021), .Q(state_1_1), .Q_N(N106), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[2] (.CLK(i_clk), .D(n1020), .Q(state_1_2), .Q_N(N117), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[3] (.CLK(i_clk), .D(n1019), .Q(state_1_3), .Q_N(N128), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[4] (.CLK(i_clk), .D(n1018), .Q(state_1_4), .Q_N(N139), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[5] (.CLK(i_clk), .D(n1017), .Q(state_1_5), .Q_N(N150), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[6] (.CLK(i_clk), .D(n1016), .Q(state_1_6), .Q_N(N161), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[7] (.CLK(i_clk), .D(n1015), .Q(state_1_7), .Q_N(N172), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[8] (.CLK(i_clk), .D(n1014), .Q(state_1_8), .Q_N(N183), .RESET_B(n1340));
sg13g2_dfrbp_1 \state_1_reg[9] (.CLK(i_clk), .D(n1023), .Q(state_1_9), .Q_N(n446), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[0] (.CLK(i_clk), .D(n940), .Q(\o_un[0]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[1] (.CLK(i_clk), .D(n939), .Q(\o_un[1]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[2] (.CLK(i_clk), .D(n938), .Q(\o_un[2]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[3] (.CLK(i_clk), .D(n937), .Q(\o_un[3]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[4] (.CLK(i_clk), .D(n936), .Q(\o_un[4]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[5] (.CLK(i_clk), .D(n935), .Q(\o_un[5]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[6] (.CLK(i_clk), .D(n934), .Q(\o_un[6]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[7] (.CLK(i_clk), .D(n933), .Q(\o_un[7]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[8] (.CLK(i_clk), .D(n932), .Q(\o_un[8]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[9] (.CLK(i_clk), .D(n931), .Q(\o_un[9]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[10] (.CLK(i_clk), .D(n930), .Q(\o_un[10]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[11] (.CLK(i_clk), .D(n929), .Q(\o_un[11]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[12] (.CLK(i_clk), .D(n928), .Q(\o_un[12]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[13] (.CLK(i_clk), .D(n927), .Q(\o_un[13]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[14] (.CLK(i_clk), .D(n926), .Q(\o_un[14]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[15] (.CLK(i_clk), .D(n925), .Q(\o_un[15]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[16] (.CLK(i_clk), .D(n924), .Q(\o_un[16]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[17] (.CLK(i_clk), .D(n923), .Q(\o_un[17]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[18] (.CLK(i_clk), .D(n922), .Q(\o_un[18]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[19] (.CLK(i_clk), .D(n921), .Q(\o_un[19]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[20] (.CLK(i_clk), .D(n920), .Q(\o_un[20]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[21] (.CLK(i_clk), .D(n919), .Q(\o_un[21]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[22] (.CLK(i_clk), .D(n918), .Q(\o_un[22]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[23] (.CLK(i_clk), .D(n917), .Q(\o_un[23]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[24] (.CLK(i_clk), .D(n916), .Q(\o_un[24]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[25] (.CLK(i_clk), .D(n915), .Q(\o_un[25]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[26] (.CLK(i_clk), .D(n914), .Q(\o_un[26]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[27] (.CLK(i_clk), .D(n913), .Q(\o_un[27]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[28] (.CLK(i_clk), .D(n912), .Q(\o_un[28]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[29] (.CLK(i_clk), .D(n911), .Q(\o_un[29]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[30] (.CLK(i_clk), .D(n910), .Q(\o_un[30]), .RESET_B(n1340));
sg13g2_dfrbp_1 \un_reg[31] (.CLK(i_clk), .D(n909), .Q(\o_un[31]), .RESET_B(n1340));
sg13g2_nand2_2 C70 (.A(n1341), .B(\i_wb_adr[3]), .Y(N48));
sg13g2_nand2_2 C74 (.A(\i_wb_adr[4]), .B(N480), .Y(N51));
sg13g2_nand2_2 C993 (.A(n410), .B(n445), .Y(N103));
sg13g2_nand2_2 C1023 (.A(N106), .B(N95), .Y(N133));
sg13g2_nand2_2 C1025 (.A(n402), .B(n421), .Y(N135));
sg13g2_nand2_2 C1034 (.A(N106), .B(N95), .Y(N144));
sg13g2_nand2_2 C1037 (.A(n410), .B(n429), .Y(N147));
sg13g2_nand2_2 C1078 (.A(N106), .B(N95), .Y(N188));
sg13g2_nand2_2 C1080 (.A(n1298), .B(n456), .Y(N190));
sg13g2_nand2_2 C1081 (.A(n451), .B(n452), .Y(N191));
sg13g2_nand2_2 C1089 (.A(N106), .B(N95), .Y(N199));
sg13g2_nand2_2 C1092 (.A(n457), .B(n445), .Y(N202));
sg13g2_nand2_2 C2587 (.A(N474), .B(mr_index_1), .Y(N478));
sg13g2_nand2_2 C2736 (.A(N522), .B(N532), .Y(n40));
sg13g2_nand2_2 C2777 (.A(N541), .B(adr_check), .Y(n36));
sg13g2_nand2_2 C2778 (.A(N540), .B(n1525), .Y(n549));
sg13g2_nand2_2 C2779 (.A(wack), .B(n1341), .Y(n550));
sg13g2_nand2_2 C2782 (.A(N542), .B(adr_check), .Y(n35));
sg13g2_nand2_2 C2783 (.A(wack), .B(N521), .Y(n551));
sg13g2_nand2_2 C2802 (.A(p_15), .B(a_15), .Y(n557));
sg13g2_nand2_2 C2805 (.A(N550), .B(N551), .Y(n559));
sg13g2_nand2_2 C2808 (.A(n560), .B(n562), .Y(\of_addition[1]));
sg13g2_nand2_2 C2809 (.A(N554), .B(n207), .Y(n560));
sg13g2_nand2_2 C2813 (.A(N557), .B(N558), .Y(n563));
sg13g2_nand2_2 C2942 (.A(re), .B(N532), .Y(n569));
sg13g2_nand2_2 C2944 (.A(re), .B(N531), .Y(n570));
sg13g2_dfrbp_1 cout_reg (.CLK(i_clk), .D(n1013), .Q(cout), .RESET_B(n1340));
sg13g2_inv_2 I_22 (.A(N39), .Y(N40));
sg13g2_dfrbp_1 rla_reg (.CLK(i_clk), .D(n1011), .Q(rl_5), .RESET_B(n1340));
sg13g2_dfrbp_1 rlb_reg (.CLK(i_clk), .D(n1009), .Q(rl_6), .Q_N(o_valid), .RESET_B(n1340));
sg13g2_dfrbp_1 RS_reg (.CLK(i_clk), .D(N81), .Q(RS), .RESET_B(n1340));
sg13g2_dfrbp_1 start_reg (.CLK(i_clk), .D(n1012), .Q(start), .RESET_B(n1340));
sg13g2_dfrbp_1 state_0_reg (.CLK(i_clk), .D(n1104), .Q(state_0), .RESET_B(n1340));
sg13g2_tielo U1 (.L_LO(n651));
sg13g2_nand3b_1 U2 (.A_N(state_1_1), .B(n18), .C(N95), .Y(n1));
sg13g2_o21ai_1 U3 (.A1(n1), .A2(n160), .B1(n2), .Y(n19));
sg13g2_nand2_2 U4 (.A(\err[1][15]), .B(n1), .Y(n2));
sg13g2_o21ai_1 U5 (.A1(n1), .A2(n164), .B1(n3), .Y(n20));
sg13g2_nand2_2 U6 (.A(\err[1][14]), .B(n1), .Y(n3));
sg13g2_o21ai_1 U7 (.A1(n1), .A2(n168), .B1(n4), .Y(n21));
sg13g2_nand2_2 U8 (.A(\err[1][13]), .B(n1), .Y(n4));
sg13g2_o21ai_1 U9 (.A1(n1), .A2(n172), .B1(n5), .Y(n22));
sg13g2_nand2_2 U10 (.A(\err[1][12]), .B(n1), .Y(n5));
sg13g2_o21ai_1 U11 (.A1(n1), .A2(n176), .B1(n6), .Y(n23));
sg13g2_nand2_2 U12 (.A(\err[1][11]), .B(n1), .Y(n6));
sg13g2_o21ai_1 U13 (.A1(n1), .A2(n180), .B1(n7), .Y(n24));
sg13g2_nand2_2 U14 (.A(\err[1][10]), .B(n1), .Y(n7));
sg13g2_o21ai_1 U15 (.A1(n1), .A2(n124), .B1(n8), .Y(n25));
sg13g2_nand2_2 U16 (.A(\err[1][9]), .B(n1), .Y(n8));
sg13g2_o21ai_1 U17 (.A1(n1), .A2(n128), .B1(n9), .Y(n26));
sg13g2_nand2_2 U18 (.A(\err[1][8]), .B(n1), .Y(n9));
sg13g2_o21ai_1 U19 (.A1(n1), .A2(n132), .B1(n10), .Y(n27));
sg13g2_nand2_2 U20 (.A(\err[1][7]), .B(n1), .Y(n10));
sg13g2_o21ai_1 U21 (.A1(n1), .A2(n136), .B1(n11), .Y(n28));
sg13g2_nand2_2 U22 (.A(\err[1][6]), .B(n1), .Y(n11));
sg13g2_o21ai_1 U23 (.A1(n1), .A2(n140), .B1(n12), .Y(n29));
sg13g2_nand2_2 U24 (.A(\err[1][5]), .B(n1), .Y(n12));
sg13g2_o21ai_1 U25 (.A1(n1), .A2(n144), .B1(n13), .Y(n30));
sg13g2_nand2_2 U26 (.A(\err[1][4]), .B(n1), .Y(n13));
sg13g2_o21ai_1 U27 (.A1(n1), .A2(n148), .B1(n14), .Y(n31));
sg13g2_nand2_2 U28 (.A(\err[1][3]), .B(n1), .Y(n14));
sg13g2_o21ai_1 U29 (.A1(n1), .A2(n152), .B1(n15), .Y(n32));
sg13g2_nand2_2 U30 (.A(\err[1][2]), .B(n1), .Y(n15));
sg13g2_o21ai_1 U31 (.A1(n1), .A2(n156), .B1(n16), .Y(n33));
sg13g2_nand2_2 U32 (.A(\err[1][1]), .B(n1), .Y(n16));
sg13g2_o21ai_1 U33 (.A1(n1), .A2(n184), .B1(n17), .Y(n34));
sg13g2_nand2_2 U34 (.A(\err[1][0]), .B(n1), .Y(n17));
sg13g2_inv_1 U35 (.A(N360), .Y(net9474));
sg13g2_inv_1 U36 (.A(n397), .Y(n376));
sg13g2_inv_1 U37 (.A(n391), .Y(n381));
sg13g2_inv_2 U38 (.A(n42), .Y(\o_wb_data[9]));
sg13g2_nand2_2 U39 (.A(N532), .B(N458), .Y(n42));
sg13g2_inv_2 U40 (.A(n43), .Y(\o_wb_data[8]));
sg13g2_nand2_2 U41 (.A(N459), .B(N532), .Y(n43));
sg13g2_inv_2 U42 (.A(n44), .Y(\o_wb_data[7]));
sg13g2_nand2_2 U43 (.A(N460), .B(N532), .Y(n44));
sg13g2_inv_2 U44 (.A(n45), .Y(\o_wb_data[6]));
sg13g2_nand2_2 U45 (.A(N461), .B(N532), .Y(n45));
sg13g2_inv_2 U46 (.A(n46), .Y(\o_wb_data[5]));
sg13g2_nand2_2 U47 (.A(N462), .B(N532), .Y(n46));
sg13g2_inv_2 U48 (.A(n47), .Y(\o_wb_data[4]));
sg13g2_nand2_2 U49 (.A(N463), .B(N532), .Y(n47));
sg13g2_inv_2 U50 (.A(n48), .Y(\o_wb_data[3]));
sg13g2_nand2_2 U51 (.A(N464), .B(N532), .Y(n48));
sg13g2_inv_2 U52 (.A(n49), .Y(\o_wb_data[31]));
sg13g2_nand2_2 U53 (.A(N436), .B(N532), .Y(n49));
sg13g2_inv_2 U54 (.A(n50), .Y(\o_wb_data[30]));
sg13g2_nand2_2 U55 (.A(N437), .B(N532), .Y(n50));
sg13g2_inv_2 U56 (.A(n51), .Y(\o_wb_data[2]));
sg13g2_nand2_2 U57 (.A(N465), .B(N532), .Y(n51));
sg13g2_inv_2 U58 (.A(n52), .Y(\o_wb_data[29]));
sg13g2_nand2_2 U59 (.A(N438), .B(N532), .Y(n52));
sg13g2_nand3b_1 U60 (.A_N(N266), .B(net9474), .C(n1), .Y(N255));
sg13g2_inv_2 U61 (.A(n53), .Y(\o_wb_data[28]));
sg13g2_nand2_2 U62 (.A(N439), .B(N532), .Y(n53));
sg13g2_inv_2 U63 (.A(n54), .Y(\o_wb_data[27]));
sg13g2_nand2_2 U64 (.A(N440), .B(N532), .Y(n54));
sg13g2_inv_2 U65 (.A(n55), .Y(\o_wb_data[26]));
sg13g2_nand2_2 U66 (.A(N441), .B(N532), .Y(n55));
sg13g2_inv_2 U67 (.A(n56), .Y(\o_wb_data[25]));
sg13g2_nand2_2 U68 (.A(N442), .B(N532), .Y(n56));
sg13g2_inv_2 U69 (.A(n57), .Y(\o_wb_data[24]));
sg13g2_nand2_2 U70 (.A(N443), .B(N532), .Y(n57));
sg13g2_inv_2 U71 (.A(n58), .Y(\o_wb_data[23]));
sg13g2_nand2_2 U72 (.A(N444), .B(N532), .Y(n58));
sg13g2_inv_2 U73 (.A(n59), .Y(\o_wb_data[22]));
sg13g2_nand2_2 U74 (.A(N445), .B(N532), .Y(n59));
sg13g2_inv_2 U75 (.A(n60), .Y(\o_wb_data[21]));
sg13g2_nand2_2 U76 (.A(N446), .B(N532), .Y(n60));
sg13g2_inv_2 U77 (.A(n61), .Y(\o_wb_data[20]));
sg13g2_nand2_2 U78 (.A(N447), .B(N532), .Y(n61));
sg13g2_inv_2 U79 (.A(n62), .Y(\o_wb_data[1]));
sg13g2_nand2_2 U80 (.A(N466), .B(N532), .Y(n62));
sg13g2_inv_2 U81 (.A(n63), .Y(\o_wb_data[19]));
sg13g2_nand2_2 U82 (.A(N448), .B(N532), .Y(n63));
sg13g2_inv_2 U83 (.A(n64), .Y(\o_wb_data[18]));
sg13g2_nand2_2 U84 (.A(N449), .B(N532), .Y(n64));
sg13g2_inv_2 U85 (.A(n65), .Y(\o_wb_data[17]));
sg13g2_nand2_2 U86 (.A(N450), .B(N532), .Y(n65));
sg13g2_inv_2 U87 (.A(n66), .Y(\o_wb_data[16]));
sg13g2_nand2_2 U88 (.A(N451), .B(N532), .Y(n66));
sg13g2_inv_2 U89 (.A(n67), .Y(\o_wb_data[15]));
sg13g2_nand2_2 U90 (.A(N452), .B(N532), .Y(n67));
sg13g2_inv_2 U91 (.A(n68), .Y(\o_wb_data[14]));
sg13g2_nand2_2 U92 (.A(N453), .B(N532), .Y(n68));
sg13g2_inv_2 U93 (.A(n69), .Y(\o_wb_data[13]));
sg13g2_nand2_2 U94 (.A(N454), .B(N532), .Y(n69));
sg13g2_inv_2 U95 (.A(n70), .Y(\o_wb_data[12]));
sg13g2_nand2_2 U96 (.A(N455), .B(N532), .Y(n70));
sg13g2_inv_2 U97 (.A(n71), .Y(\o_wb_data[11]));
sg13g2_nand2_2 U98 (.A(N456), .B(N532), .Y(n71));
sg13g2_inv_2 U99 (.A(n72), .Y(\o_wb_data[10]));
sg13g2_nand2_2 U100 (.A(N457), .B(N532), .Y(n72));
sg13g2_inv_2 U101 (.A(n73), .Y(\o_wb_data[0]));
sg13g2_nand2_2 U102 (.A(N467), .B(N532), .Y(n73));
sg13g2_o21ai_1 U103 (.A1(n388), .A2(n35), .B1(n37), .Y(N266));
sg13g2_nand2_2 U104 (.A(ki_9), .B(N91), .Y(n77));
sg13g2_nand2_2 U105 (.A(kpd_9), .B(N476), .Y(n76));
sg13g2_o21ai_1 U106 (.A1(n39), .A2(n41), .B1(n74), .Y(n652));
sg13g2_nand3_1 U107 (.A(n311), .B(n75), .C(n310), .Y(n293));
sg13g2_nand2_2 U108 (.A(ki_8), .B(N91), .Y(n80));
sg13g2_nand2_2 U109 (.A(kpd_8), .B(N476), .Y(n79));
sg13g2_nand3_1 U110 (.A(n284), .B(n78), .C(n283), .Y(N394));
sg13g2_nand3_1 U111 (.A(n257), .B(n81), .C(n256), .Y(N403));
sg13g2_nand2_2 U112 (.A(ki_7), .B(N91), .Y(n83));
sg13g2_nand2_2 U113 (.A(kpd_7), .B(N476), .Y(n82));
sg13g2_nand2_1 U114 (.A(n84), .B(n216), .Y(N421));
sg13g2_nand2_1 U115 (.A(n87), .B(n224), .Y(N417));
sg13g2_nand2_2 U116 (.A(ki_6), .B(N91), .Y(n86));
sg13g2_nand2_2 U117 (.A(kpd_6), .B(N476), .Y(n85));
sg13g2_nand3_1 U118 (.A(n245), .B(n90), .C(n244), .Y(N407));
sg13g2_nand2_1 U119 (.A(n93), .B(n236), .Y(N411));
sg13g2_nand2_2 U120 (.A(ki_5), .B(N91), .Y(n89));
sg13g2_nand2_2 U121 (.A(kpd_5), .B(N476), .Y(n88));
sg13g2_nand3_1 U122 (.A(n263), .B(n96), .C(n262), .Y(N401));
sg13g2_nand2_1 U123 (.A(n99), .B(n228), .Y(N415));
sg13g2_nand2_2 U124 (.A(ki_4), .B(N91), .Y(n92));
sg13g2_nand2_2 U125 (.A(kpd_4), .B(N476), .Y(n91));
sg13g2_nand2_1 U126 (.A(n102), .B(n212), .Y(N423));
sg13g2_nand3_1 U127 (.A(n254), .B(n105), .C(n253), .Y(N404));
sg13g2_nand2_2 U128 (.A(ki_3), .B(N91), .Y(n95));
sg13g2_nand2_2 U129 (.A(kpd_3), .B(N476), .Y(n94));
sg13g2_nand2_1 U130 (.A(n108), .B(n240), .Y(N409));
sg13g2_nand3_1 U131 (.A(n260), .B(n111), .C(n259), .Y(N402));
sg13g2_nand2_2 U132 (.A(ki_2), .B(N91), .Y(n98));
sg13g2_nand2_2 U133 (.A(kpd_2), .B(N476), .Y(n97));
sg13g2_nand2_1 U134 (.A(n114), .B(n230), .Y(N414));
sg13g2_nand2_1 U135 (.A(n117), .B(n232), .Y(N413));
sg13g2_nand2_2 U136 (.A(ki_1), .B(N91), .Y(n101));
sg13g2_nand2_2 U137 (.A(kpd_1), .B(N476), .Y(n100));
sg13g2_nand3_1 U138 (.A(n281), .B(n120), .C(n280), .Y(N395));
sg13g2_nand3_1 U139 (.A(n275), .B(n188), .C(n274), .Y(N397));
sg13g2_nand2_2 U140 (.A(ki_15), .B(N91), .Y(n104));
sg13g2_nand2_2 U141 (.A(kpd_15), .B(N476), .Y(n103));
sg13g2_a21oi_1 U142 (.A1(n189), .A2(n568), .B1(n1276), .Y(o_wb_ack));
sg13g2_nand3_1 U143 (.A(n272), .B(n191), .C(n271), .Y(N398));
sg13g2_nand2_2 U144 (.A(ki_14), .B(N91), .Y(n107));
sg13g2_nand2_2 U145 (.A(kpd_14), .B(N476), .Y(n106));
sg13g2_nand3_1 U146 (.A(n269), .B(n192), .C(n268), .Y(N399));
sg13g2_nand3_1 U147 (.A(n266), .B(n193), .C(n265), .Y(N400));
sg13g2_nand2_2 U148 (.A(ki_13), .B(N91), .Y(n110));
sg13g2_nand2_2 U149 (.A(kpd_13), .B(N476), .Y(n109));
sg13g2_nand3_1 U150 (.A(n248), .B(n195), .C(n247), .Y(N406));
sg13g2_nand3_1 U151 (.A(n251), .B(n197), .C(n250), .Y(N405));
sg13g2_nand2_2 U152 (.A(ki_12), .B(N91), .Y(n113));
sg13g2_nand2_2 U153 (.A(kpd_12), .B(N476), .Y(n112));
sg13g2_nand2_1 U154 (.A(n198), .B(n220), .Y(N419));
sg13g2_nand3_1 U155 (.A(n278), .B(n201), .C(n277), .Y(N396));
sg13g2_nand2_2 U156 (.A(ki_11), .B(N91), .Y(n116));
sg13g2_nand2_2 U157 (.A(kpd_11), .B(N476), .Y(n115));
sg13g2_nand2_1 U158 (.A(n202), .B(n241), .Y(N408));
sg13g2_nand2_1 U159 (.A(n203), .B(n238), .Y(N410));
sg13g2_nand2_2 U160 (.A(ki_10), .B(N91), .Y(n119));
sg13g2_nand2_2 U161 (.A(kpd_10), .B(N476), .Y(n118));
sg13g2_nand2_1 U162 (.A(n209), .B(n234), .Y(N412));
sg13g2_nand2_1 U163 (.A(n298), .B(n226), .Y(N416));
sg13g2_nand2_2 U164 (.A(ki_0), .B(N91), .Y(n122));
sg13g2_nand2_2 U165 (.A(kpd_0), .B(N476), .Y(n121));
sg13g2_nand2_1 U166 (.A(n301), .B(n222), .Y(N418));
sg13g2_nand2_1 U167 (.A(n382), .B(n218), .Y(N420));
sg13g2_o21ai_1 U168 (.A1(n123), .A2(n124), .B1(n125), .Y(md_9));
sg13g2_a21oi_2 U169 (.A1(\err[1][9]), .A2(N470), .B1(n126), .Y(n125));
sg13g2_inv_2 U170 (.A(n127), .Y(n126));
sg13g2_nand2_2 U171 (.A(N473), .B(\err[0][9]), .Y(n127));
sg13g2_o21ai_1 U172 (.A1(n123), .A2(n128), .B1(n129), .Y(md_8));
sg13g2_a21oi_2 U173 (.A1(\err[1][8]), .A2(N470), .B1(n130), .Y(n129));
sg13g2_inv_2 U174 (.A(n131), .Y(n130));
sg13g2_nand2_2 U175 (.A(N473), .B(\err[0][8]), .Y(n131));
sg13g2_o21ai_1 U176 (.A1(n123), .A2(n132), .B1(n133), .Y(md_7));
sg13g2_a21oi_2 U177 (.A1(\err[1][7]), .A2(N470), .B1(n134), .Y(n133));
sg13g2_inv_2 U178 (.A(n135), .Y(n134));
sg13g2_nand2_2 U179 (.A(N473), .B(\err[0][7]), .Y(n135));
sg13g2_o21ai_1 U180 (.A1(n123), .A2(n136), .B1(n137), .Y(md_6));
sg13g2_a21oi_2 U181 (.A1(\err[1][6]), .A2(N470), .B1(n138), .Y(n137));
sg13g2_inv_2 U182 (.A(n139), .Y(n138));
sg13g2_nand2_2 U183 (.A(N473), .B(\err[0][6]), .Y(n139));
sg13g2_o21ai_1 U184 (.A1(n123), .A2(n140), .B1(n141), .Y(md_5));
sg13g2_a21oi_2 U185 (.A1(\err[1][5]), .A2(N470), .B1(n142), .Y(n141));
sg13g2_inv_2 U186 (.A(n143), .Y(n142));
sg13g2_nand2_2 U187 (.A(N473), .B(\err[0][5]), .Y(n143));
sg13g2_o21ai_1 U188 (.A1(n123), .A2(n144), .B1(n145), .Y(md_4));
sg13g2_a21oi_2 U189 (.A1(\err[1][4]), .A2(N470), .B1(n146), .Y(n145));
sg13g2_inv_2 U190 (.A(n147), .Y(n146));
sg13g2_nand2_2 U191 (.A(N473), .B(\err[0][4]), .Y(n147));
sg13g2_o21ai_1 U192 (.A1(n123), .A2(n148), .B1(n149), .Y(md_3));
sg13g2_a21oi_2 U193 (.A1(\err[1][3]), .A2(N470), .B1(n150), .Y(n149));
sg13g2_inv_2 U194 (.A(n151), .Y(n150));
sg13g2_nand2_2 U195 (.A(N473), .B(\err[0][3]), .Y(n151));
sg13g2_o21ai_1 U196 (.A1(n123), .A2(n152), .B1(n153), .Y(md_2));
sg13g2_a21oi_2 U197 (.A1(\err[1][2]), .A2(N470), .B1(n154), .Y(n153));
sg13g2_inv_2 U198 (.A(n155), .Y(n154));
sg13g2_nand2_2 U199 (.A(N473), .B(\err[0][2]), .Y(n155));
sg13g2_o21ai_1 U200 (.A1(n123), .A2(n156), .B1(n157), .Y(md_1));
sg13g2_a21oi_2 U201 (.A1(\err[1][1]), .A2(N470), .B1(n158), .Y(n157));
sg13g2_inv_2 U202 (.A(n159), .Y(n158));
sg13g2_nand2_2 U203 (.A(N473), .B(\err[0][1]), .Y(n159));
sg13g2_nand2_1 U204 (.A(n383), .B(n214), .Y(N422));
sg13g2_a21oi_2 U205 (.A1(\err[1][15]), .A2(N470), .B1(n162), .Y(n161));
sg13g2_inv_2 U206 (.A(n163), .Y(n162));
sg13g2_nand2_2 U207 (.A(N473), .B(\err[0][15]), .Y(n163));
sg13g2_o21ai_1 U208 (.A1(n123), .A2(n164), .B1(n165), .Y(md_14));
sg13g2_a21oi_2 U209 (.A1(\err[1][14]), .A2(N470), .B1(n166), .Y(n165));
sg13g2_inv_2 U210 (.A(n167), .Y(n166));
sg13g2_nand2_2 U211 (.A(N473), .B(\err[0][14]), .Y(n167));
sg13g2_o21ai_1 U212 (.A1(n123), .A2(n168), .B1(n169), .Y(md_13));
sg13g2_a21oi_2 U213 (.A1(\err[1][13]), .A2(N470), .B1(n170), .Y(n169));
sg13g2_inv_2 U214 (.A(n171), .Y(n170));
sg13g2_nand2_2 U215 (.A(N473), .B(\err[0][13]), .Y(n171));
sg13g2_nand2_1 U216 (.A(n386), .B(n210), .Y(N424));
sg13g2_a21oi_2 U217 (.A1(\err[1][12]), .A2(N470), .B1(n174), .Y(n173));
sg13g2_inv_2 U218 (.A(n175), .Y(n174));
sg13g2_nand2_2 U219 (.A(N473), .B(\err[0][12]), .Y(n175));
sg13g2_o21ai_1 U220 (.A1(n123), .A2(n176), .B1(n177), .Y(md_11));
sg13g2_a21oi_2 U221 (.A1(\err[1][11]), .A2(N470), .B1(n178), .Y(n177));
sg13g2_inv_2 U222 (.A(n179), .Y(n178));
sg13g2_nand2_2 U223 (.A(N473), .B(\err[0][11]), .Y(n179));
sg13g2_o21ai_1 U224 (.A1(n123), .A2(n180), .B1(n181), .Y(md_10));
sg13g2_a21oi_2 U225 (.A1(\err[1][10]), .A2(N470), .B1(n182), .Y(n181));
sg13g2_inv_2 U226 (.A(n183), .Y(n182));
sg13g2_nand2_2 U227 (.A(N473), .B(\err[0][10]), .Y(n183));
sg13g2_o21ai_1 U228 (.A1(n123), .A2(n184), .B1(n185), .Y(md_0));
sg13g2_a21oi_2 U229 (.A1(\err[1][0]), .A2(N470), .B1(n186), .Y(n185));
sg13g2_inv_2 U230 (.A(n187), .Y(n186));
sg13g2_nand2_2 U231 (.A(N473), .B(\err[0][0]), .Y(n187));
sg13g2_nand3_1 U232 (.A(n77), .B(n387), .C(n76), .Y(mr_9));
sg13g2_nand3_1 U233 (.A(n80), .B(n394), .C(n79), .Y(mr_8));
sg13g2_nand3_1 U234 (.A(n83), .B(n400), .C(n82), .Y(mr_7));
sg13g2_nand3_1 U235 (.A(n86), .B(n401), .C(n85), .Y(mr_6));
sg13g2_nand3_1 U236 (.A(n89), .B(n403), .C(n88), .Y(mr_5));
sg13g2_nand3_1 U237 (.A(n92), .B(n404), .C(n91), .Y(mr_4));
sg13g2_nand3_1 U238 (.A(n95), .B(n405), .C(n94), .Y(mr_3));
sg13g2_nand3_1 U239 (.A(n98), .B(n406), .C(n97), .Y(mr_2));
sg13g2_nand3_1 U240 (.A(n101), .B(n407), .C(n100), .Y(mr_1));
sg13g2_nand3_1 U241 (.A(n104), .B(n408), .C(n103), .Y(mr_15));
sg13g2_nand3_1 U242 (.A(n107), .B(n409), .C(n106), .Y(mr_14));
sg13g2_nand3_1 U243 (.A(n110), .B(n411), .C(n109), .Y(mr_13));
sg13g2_nand3_1 U244 (.A(n113), .B(n412), .C(n112), .Y(mr_12));
sg13g2_inv_2 U245 (.A(n196), .Y(n190));
sg13g2_nand3_1 U246 (.A(N40), .B(adr_check), .C(state_0), .Y(n196));
sg13g2_nand3_1 U247 (.A(n116), .B(n414), .C(n115), .Y(mr_11));
sg13g2_nand3_1 U248 (.A(n119), .B(n417), .C(n118), .Y(mr_10));
sg13g2_nand3_1 U249 (.A(n122), .B(n418), .C(n121), .Y(mr_0));
sg13g2_o21ai_1 U250 (.A1(state_0), .A2(n38), .B1(n194), .Y(N79));
sg13g2_o21ai_1 U251 (.A1(N40), .A2(n40), .B1(state_0), .Y(n194));
sg13g2_nor2b_1 U252 (.A(state_1_1), .B_N(n18), .Y(n419));
sg13g2_inv_2 U253 (.A(N51), .Y(n199));
sg13g2_nor3_1 U254 (.A(n419), .B(N360), .C(N266), .Y(n39));
sg13g2_nor2_1 U255 (.A(n391), .B(n397), .Y(n41));
sg13g2_inv_2 U256 (.A(N48), .Y(n200));
sg13g2_nor2_1 U257 (.A(n391), .B(N268), .Y(n37));
sg13g2_and2_1 U258 (.A(n570), .B(N537), .X(n189));
sg13g2_a21oi_1 U259 (.A1(n1291), .A2(sum_31), .B1(n242), .Y(n386));
sg13g2_a21oi_1 U260 (.A1(n1291), .A2(sum_30), .B1(n242), .Y(n102));
sg13g2_inv_2 U261 (.A(n205), .Y(N427));
sg13g2_nand2_2 U262 (.A(n204), .B(n206), .Y(N426));
sg13g2_a21oi_1 U263 (.A1(n1291), .A2(sum_29), .B1(n242), .Y(n383));
sg13g2_a21oi_1 U264 (.A1(n1291), .A2(sum_28), .B1(n242), .Y(n84));
sg13g2_a21oi_1 U265 (.A1(n1291), .A2(sum_27), .B1(n242), .Y(n382));
sg13g2_a21oi_1 U266 (.A1(n1291), .A2(sum_26), .B1(n242), .Y(n198));
sg13g2_a21oi_1 U267 (.A1(n1291), .A2(sum_25), .B1(n242), .Y(n301));
sg13g2_a21oi_2 U268 (.A1(sigma_29), .A2(N263), .B1(N333), .Y(n214));
sg13g2_a21oi_1 U269 (.A1(n1291), .A2(sum_24), .B1(n242), .Y(n87));
sg13g2_a21oi_1 U270 (.A1(n1291), .A2(sum_23), .B1(n242), .Y(n298));
sg13g2_a21oi_1 U271 (.A1(n1291), .A2(sum_22), .B1(n242), .Y(n99));
sg13g2_a21oi_1 U272 (.A1(n1291), .A2(sum_21), .B1(n242), .Y(n114));
sg13g2_a21oi_1 U273 (.A1(n1291), .A2(sum_20), .B1(n242), .Y(n117));
sg13g2_a21oi_1 U274 (.A1(n1291), .A2(sum_19), .B1(n242), .Y(n209));
sg13g2_a21oi_1 U275 (.A1(n1291), .A2(sum_18), .B1(n242), .Y(n93));
sg13g2_a21oi_1 U276 (.A1(n1291), .A2(sum_17), .B1(n242), .Y(n203));
sg13g2_a21oi_1 U277 (.A1(n1291), .A2(sum_16), .B1(n242), .Y(n108));
sg13g2_a21oi_1 U278 (.A1(n1291), .A2(sum_15), .B1(n242), .Y(n202));
sg13g2_inv_1 U279 (.A(N478), .Y(n420));
sg13g2_or3_1 U280 (.A(N95), .B(N360), .C(N266), .X(n74));
sg13g2_nand2_1 U281 (.A(n395), .B(n422), .Y(n75));
sg13g2_nand2_1 U282 (.A(kd_9), .B(n420), .Y(n387));
sg13g2_nand2_1 U283 (.A(kd_8), .B(n420), .Y(n394));
sg13g2_a21oi_2 U284 (.A1(sigma_21), .A2(N263), .B1(N325), .Y(n230));
sg13g2_nand2_1 U285 (.A(kd_7), .B(n420), .Y(n400));
sg13g2_a21oi_2 U286 (.A1(sigma_20), .A2(N263), .B1(N324), .Y(n232));
sg13g2_nand2_1 U287 (.A(kd_6), .B(n420), .Y(n401));
sg13g2_a21oi_2 U288 (.A1(sigma_19), .A2(N263), .B1(N323), .Y(n234));
sg13g2_nand2_1 U289 (.A(kd_5), .B(n420), .Y(n403));
sg13g2_nand2_1 U290 (.A(kd_4), .B(n420), .Y(n404));
sg13g2_nand2_1 U291 (.A(kd_3), .B(n420), .Y(n405));
sg13g2_a21oi_2 U292 (.A1(sigma_17), .A2(N263), .B1(N321), .Y(n238));
sg13g2_nand2_1 U293 (.A(kd_2), .B(n420), .Y(n406));
sg13g2_nand2_1 U294 (.A(kd_1), .B(n420), .Y(n407));
sg13g2_nand2_1 U295 (.A(kd_15), .B(n420), .Y(n408));
sg13g2_a21oi_2 U296 (.A1(sigma_15), .A2(N263), .B1(N319), .Y(n241));
sg13g2_nand2_1 U297 (.A(kd_14), .B(n420), .Y(n409));
sg13g2_nand2_1 U298 (.A(kd_13), .B(n420), .Y(n411));
sg13g2_nand2_2 U299 (.A(n398), .B(kd_15), .Y(n243));
sg13g2_nand2_1 U300 (.A(kd_12), .B(n420), .Y(n412));
sg13g2_nand2_1 U301 (.A(kd_11), .B(n420), .Y(n414));
sg13g2_nand2_1 U302 (.A(kd_10), .B(n420), .Y(n417));
sg13g2_nand2_1 U303 (.A(kd_0), .B(n420), .Y(n418));
sg13g2_nand2_1 U304 (.A(n396), .B(n427), .Y(n90));
sg13g2_a21oi_2 U305 (.A1(sigma_13), .A2(N263), .B1(n249), .Y(n248));
sg13g2_nor2_2 U306 (.A(n168), .B(n208), .Y(n249));
sg13g2_a21oi_2 U307 (.A1(n398), .A2(kd_13), .B1(N317), .Y(n247));
sg13g2_nand2_1 U308 (.A(n396), .B(n440), .Y(n195));
sg13g2_a21oi_2 U309 (.A1(sigma_12), .A2(N263), .B1(n252), .Y(n251));
sg13g2_nand2_1 U310 (.A(n396), .B(n441), .Y(n197));
sg13g2_nand2_1 U311 (.A(n396), .B(n433), .Y(n105));
sg13g2_nand2_1 U312 (.A(n396), .B(n425), .Y(n81));
sg13g2_a21oi_2 U313 (.A1(sigma_11), .A2(N263), .B1(n255), .Y(n254));
sg13g2_nor2_2 U314 (.A(n176), .B(n208), .Y(n255));
sg13g2_a21oi_2 U315 (.A1(n398), .A2(kd_11), .B1(N315), .Y(n253));
sg13g2_nand2_1 U316 (.A(n396), .B(n434), .Y(n111));
sg13g2_a21oi_2 U317 (.A1(sigma_10), .A2(N263), .B1(n258), .Y(n257));
sg13g2_nor2_2 U318 (.A(n180), .B(n208), .Y(n258));
sg13g2_a21oi_2 U319 (.A1(n398), .A2(kd_10), .B1(N314), .Y(n256));
sg13g2_nand2_1 U320 (.A(n396), .B(n428), .Y(n96));
sg13g2_a21oi_2 U321 (.A1(sigma_9), .A2(N263), .B1(n261), .Y(n260));
sg13g2_nor2_2 U322 (.A(n124), .B(n208), .Y(n261));
sg13g2_a21oi_2 U323 (.A1(n398), .A2(kd_9), .B1(N313), .Y(n259));
sg13g2_nand2_1 U324 (.A(n396), .B(n439), .Y(n193));
sg13g2_a21oi_2 U325 (.A1(sigma_8), .A2(N263), .B1(n264), .Y(n263));
sg13g2_nor2_2 U326 (.A(n128), .B(n208), .Y(n264));
sg13g2_a21oi_2 U327 (.A1(n398), .A2(kd_8), .B1(N312), .Y(n262));
sg13g2_nand2_1 U328 (.A(n396), .B(n438), .Y(n192));
sg13g2_a21oi_2 U329 (.A1(sigma_7), .A2(N263), .B1(n267), .Y(n266));
sg13g2_nor2_2 U330 (.A(n132), .B(n208), .Y(n267));
sg13g2_a21oi_2 U331 (.A1(n398), .A2(kd_7), .B1(N311), .Y(n265));
sg13g2_nand2_1 U332 (.A(n396), .B(n437), .Y(n191));
sg13g2_a21oi_2 U333 (.A1(sigma_6), .A2(N263), .B1(n270), .Y(n269));
sg13g2_nor2_2 U334 (.A(n136), .B(n208), .Y(n270));
sg13g2_a21oi_2 U335 (.A1(n398), .A2(kd_6), .B1(N310), .Y(n268));
sg13g2_nand2_1 U336 (.A(n396), .B(n436), .Y(n188));
sg13g2_a21oi_2 U337 (.A1(sigma_5), .A2(N263), .B1(n273), .Y(n272));
sg13g2_nor2_2 U338 (.A(n140), .B(n208), .Y(n273));
sg13g2_a21oi_2 U339 (.A1(n398), .A2(kd_5), .B1(N309), .Y(n271));
sg13g2_nand2_1 U340 (.A(n396), .B(n442), .Y(n201));
sg13g2_a21oi_2 U341 (.A1(sigma_4), .A2(N263), .B1(n276), .Y(n275));
sg13g2_nor2_2 U342 (.A(n144), .B(n208), .Y(n276));
sg13g2_a21oi_2 U343 (.A1(n398), .A2(kd_4), .B1(N308), .Y(n274));
sg13g2_nand2_1 U344 (.A(n396), .B(n435), .Y(n120));
sg13g2_a21oi_2 U345 (.A1(sigma_3), .A2(N263), .B1(n279), .Y(n278));
sg13g2_nor2_2 U346 (.A(n148), .B(n208), .Y(n279));
sg13g2_a21oi_2 U347 (.A1(n398), .A2(kd_3), .B1(N307), .Y(n277));
sg13g2_nand2_1 U348 (.A(n396), .B(n424), .Y(n78));
sg13g2_a21oi_2 U349 (.A1(sigma_2), .A2(N263), .B1(n282), .Y(n281));
sg13g2_nor2_2 U350 (.A(n152), .B(n208), .Y(n282));
sg13g2_a21oi_2 U351 (.A1(n398), .A2(kd_2), .B1(N306), .Y(n280));
sg13g2_inv_2 U352 (.A(n443), .Y(net9912));
sg13g2_a21oi_2 U353 (.A1(sigma_1), .A2(N263), .B1(n285), .Y(n284));
sg13g2_nor2_2 U354 (.A(n156), .B(n208), .Y(n285));
sg13g2_a21oi_2 U355 (.A1(n398), .A2(kd_1), .B1(N305), .Y(n283));
sg13g2_nand4_1 U356 (.A(n286), .B(n204), .C(n287), .D(n288), .Y(N393));
sg13g2_a21oi_2 U357 (.A1(n392), .A2(sum_0), .B1(n289), .Y(n288));
sg13g2_inv_2 U358 (.A(n447), .Y(n1305));
sg13g2_nand2_2 U359 (.A(sigma_0), .B(N263), .Y(n290));
sg13g2_inv_2 U360 (.A(n448), .Y(n1311));
sg13g2_nand2_2 U361 (.A(n398), .B(kd_0), .Y(n287));
sg13g2_inv_2 U362 (.A(N304), .Y(n286));
sg13g2_inv_2 U363 (.A(n449), .Y(n1327));
sg13g2_inv_2 U364 (.A(n450), .Y(n1300));
sg13g2_inv_2 U365 (.A(n453), .Y(n1309));
sg13g2_inv_2 U366 (.A(n454), .Y(n1325));
sg13g2_inv_2 U367 (.A(n455), .Y(n1347));
sg13g2_inv_2 U368 (.A(n458), .Y(n1350));
sg13g2_inv_2 U369 (.A(n459), .Y(N436));
sg13g2_inv_2 U370 (.A(n460), .Y(N437));
sg13g2_inv_2 U371 (.A(n461), .Y(N438));
sg13g2_inv_2 U372 (.A(n462), .Y(N439));
sg13g2_inv_2 U373 (.A(n464), .Y(N440));
sg13g2_inv_2 U374 (.A(n466), .Y(N441));
sg13g2_inv_2 U375 (.A(n299), .Y(N386));
sg13g2_a21oi_2 U376 (.A1(product_25), .A2(n292), .B1(n293), .Y(n299));
sg13g2_inv_2 U377 (.A(n467), .Y(N442));
sg13g2_inv_2 U378 (.A(n468), .Y(N443));
sg13g2_inv_2 U379 (.A(n469), .Y(N444));
sg13g2_inv_2 U380 (.A(n470), .Y(N445));
sg13g2_inv_2 U381 (.A(n473), .Y(N446));
sg13g2_inv_2 U382 (.A(n474), .Y(N447));
sg13g2_inv_2 U383 (.A(n476), .Y(N448));
sg13g2_inv_2 U384 (.A(n477), .Y(N449));
sg13g2_inv_2 U385 (.A(n478), .Y(N450));
sg13g2_inv_2 U386 (.A(n479), .Y(N451));
sg13g2_inv_2 U387 (.A(n480), .Y(N452));
sg13g2_inv_2 U388 (.A(n482), .Y(n1388));
sg13g2_inv_2 U389 (.A(n484), .Y(n1391));
sg13g2_inv_2 U390 (.A(n485), .Y(N453));
sg13g2_inv_2 U391 (.A(n307), .Y(N378));
sg13g2_a21oi_2 U392 (.A1(n292), .A2(product_17), .B1(n293), .Y(n307));
sg13g2_inv_2 U393 (.A(n486), .Y(n1397));
sg13g2_inv_2 U394 (.A(n488), .Y(n1400));
sg13g2_inv_2 U395 (.A(n309), .Y(N376));
sg13g2_a21oi_2 U396 (.A1(product_15), .A2(n292), .B1(n293), .Y(n309));
sg13g2_inv_2 U397 (.A(n490), .Y(N454));
sg13g2_nand2_2 U398 (.A(kp_15), .B(n398), .Y(n311));
sg13g2_nand2_2 U399 (.A(sp_15), .B(n396), .Y(n310));
sg13g2_inv_2 U400 (.A(n491), .Y(n1406));
sg13g2_a21oi_2 U401 (.A1(sp_14), .A2(n396), .B1(n315), .Y(n314));
sg13g2_nor2_2 U402 (.A(\err[0][14]), .B(n204), .Y(n315));
sg13g2_inv_2 U403 (.A(n492), .Y(n1409));
sg13g2_nand2_2 U404 (.A(kp_14), .B(n398), .Y(n312));
sg13g2_inv_2 U405 (.A(n494), .Y(N455));
sg13g2_a21oi_2 U406 (.A1(sp_13), .A2(n396), .B1(n319), .Y(n318));
sg13g2_nor2_2 U407 (.A(\err[0][13]), .B(n204), .Y(n319));
sg13g2_nand2_2 U408 (.A(product_13), .B(n292), .Y(n317));
sg13g2_nand2_2 U409 (.A(kp_13), .B(n398), .Y(n316));
sg13g2_inv_2 U410 (.A(n495), .Y(n1415));
sg13g2_a21oi_2 U411 (.A1(sp_12), .A2(n396), .B1(n323), .Y(n322));
sg13g2_nor2_2 U412 (.A(\err[0][12]), .B(n204), .Y(n323));
sg13g2_inv_2 U413 (.A(n496), .Y(n1418));
sg13g2_nand2_2 U414 (.A(kp_12), .B(n398), .Y(n320));
sg13g2_inv_2 U415 (.A(n497), .Y(N456));
sg13g2_a21oi_2 U416 (.A1(sp_11), .A2(n396), .B1(n327), .Y(n326));
sg13g2_nor2_2 U417 (.A(\err[0][11]), .B(n204), .Y(n327));
sg13g2_nand2_2 U418 (.A(product_11), .B(n292), .Y(n325));
sg13g2_nand2_2 U419 (.A(kp_11), .B(n398), .Y(n324));
sg13g2_inv_2 U420 (.A(n498), .Y(n1424));
sg13g2_a21oi_2 U421 (.A1(sp_10), .A2(n396), .B1(n331), .Y(n330));
sg13g2_nor2_2 U422 (.A(\err[0][10]), .B(n204), .Y(n331));
sg13g2_inv_2 U423 (.A(n500), .Y(n1427));
sg13g2_nand2_2 U424 (.A(kp_10), .B(n398), .Y(n328));
sg13g2_inv_2 U425 (.A(n502), .Y(N457));
sg13g2_a21oi_2 U426 (.A1(sp_9), .A2(n396), .B1(n335), .Y(n334));
sg13g2_nor2_2 U427 (.A(\err[0][9]), .B(n204), .Y(n335));
sg13g2_nand2_2 U428 (.A(product_9), .B(n292), .Y(n333));
sg13g2_nand2_2 U429 (.A(kp_9), .B(n398), .Y(n332));
sg13g2_inv_2 U430 (.A(n503), .Y(n1433));
sg13g2_a21oi_2 U431 (.A1(sp_8), .A2(n396), .B1(n339), .Y(n338));
sg13g2_nor2_2 U432 (.A(\err[0][8]), .B(n204), .Y(n339));
sg13g2_nand2_2 U433 (.A(product_8), .B(n292), .Y(n337));
sg13g2_nand2_2 U434 (.A(kp_8), .B(n398), .Y(n336));
sg13g2_inv_2 U435 (.A(n504), .Y(n1436));
sg13g2_a21oi_2 U436 (.A1(sp_7), .A2(n396), .B1(n343), .Y(n342));
sg13g2_nor2_2 U437 (.A(\err[0][7]), .B(n204), .Y(n343));
sg13g2_nand2_2 U438 (.A(product_7), .B(n292), .Y(n341));
sg13g2_nand2_2 U439 (.A(kp_7), .B(n398), .Y(n340));
sg13g2_inv_2 U440 (.A(n505), .Y(N458));
sg13g2_a21oi_2 U441 (.A1(sp_6), .A2(n396), .B1(n347), .Y(n346));
sg13g2_nor2_2 U442 (.A(\err[0][6]), .B(n204), .Y(n347));
sg13g2_nand2_2 U443 (.A(product_6), .B(n292), .Y(n345));
sg13g2_nand2_2 U444 (.A(kp_6), .B(n398), .Y(n344));
sg13g2_inv_2 U445 (.A(n506), .Y(n1442));
sg13g2_a21oi_2 U446 (.A1(sp_5), .A2(n396), .B1(n351), .Y(n350));
sg13g2_nor2_2 U447 (.A(\err[0][5]), .B(n204), .Y(n351));
sg13g2_nand2_2 U448 (.A(product_5), .B(n292), .Y(n349));
sg13g2_nand2_2 U449 (.A(kp_5), .B(n398), .Y(n348));
sg13g2_inv_2 U450 (.A(n509), .Y(n1445));
sg13g2_a21oi_2 U451 (.A1(sp_4), .A2(n396), .B1(n355), .Y(n354));
sg13g2_nor2_2 U452 (.A(\err[0][4]), .B(n204), .Y(n355));
sg13g2_nand2_2 U453 (.A(product_4), .B(n292), .Y(n353));
sg13g2_nand2_2 U454 (.A(kp_4), .B(n398), .Y(n352));
sg13g2_inv_2 U455 (.A(n510), .Y(N459));
sg13g2_a21oi_2 U456 (.A1(sp_3), .A2(n396), .B1(n359), .Y(n358));
sg13g2_nor2_2 U457 (.A(\err[0][3]), .B(n204), .Y(n359));
sg13g2_nand2_2 U458 (.A(product_3), .B(n292), .Y(n357));
sg13g2_nand2_2 U459 (.A(kp_3), .B(n398), .Y(n356));
sg13g2_inv_2 U460 (.A(n512), .Y(n1451));
sg13g2_a21oi_2 U461 (.A1(sp_2), .A2(n396), .B1(n363), .Y(n362));
sg13g2_nor2_2 U462 (.A(\err[0][2]), .B(n204), .Y(n363));
sg13g2_nand2_2 U463 (.A(product_2), .B(n292), .Y(n361));
sg13g2_nand2_2 U464 (.A(kp_2), .B(n398), .Y(n360));
sg13g2_inv_2 U465 (.A(n515), .Y(n1454));
sg13g2_a21oi_2 U466 (.A1(sp_1), .A2(n396), .B1(n367), .Y(n366));
sg13g2_nor2_2 U467 (.A(\err[0][1]), .B(n204), .Y(n367));
sg13g2_nand2_2 U468 (.A(product_1), .B(n292), .Y(n365));
sg13g2_nand2_2 U469 (.A(kp_1), .B(n398), .Y(n364));
sg13g2_inv_2 U470 (.A(n516), .Y(N460));
sg13g2_a21oi_2 U471 (.A1(sp_0), .A2(n396), .B1(n371), .Y(n370));
sg13g2_nor2_2 U472 (.A(\err[0][0]), .B(n204), .Y(n371));
sg13g2_nand2_2 U473 (.A(product_0), .B(n292), .Y(n369));
sg13g2_inv_2 U474 (.A(n518), .Y(n1460));
sg13g2_inv_2 U475 (.A(n519), .Y(n1463));
sg13g2_inv_2 U476 (.A(n520), .Y(N461));
sg13g2_nand2_2 U477 (.A(kp_0), .B(n398), .Y(n368));
sg13g2_nor2_2 U478 (.A(n160), .B(n204), .Y(N359));
sg13g2_nor2_2 U479 (.A(n164), .B(n204), .Y(N358));
sg13g2_nor2_2 U480 (.A(n168), .B(n204), .Y(N357));
sg13g2_nor2_2 U481 (.A(n172), .B(n204), .Y(N356));
sg13g2_nor2_2 U482 (.A(n176), .B(n204), .Y(N355));
sg13g2_nor2_2 U483 (.A(n180), .B(n204), .Y(N354));
sg13g2_nor2_2 U484 (.A(n124), .B(n204), .Y(N353));
sg13g2_nor2_2 U485 (.A(n128), .B(n204), .Y(N352));
sg13g2_nor2_2 U486 (.A(n132), .B(n204), .Y(N351));
sg13g2_nor2_2 U487 (.A(n136), .B(n204), .Y(N350));
sg13g2_nor2_2 U488 (.A(n140), .B(n204), .Y(N349));
sg13g2_nor2_2 U489 (.A(n144), .B(n204), .Y(N348));
sg13g2_nor2_2 U490 (.A(n148), .B(n204), .Y(N347));
sg13g2_nor2_2 U491 (.A(n152), .B(n204), .Y(N346));
sg13g2_nor2_2 U492 (.A(n156), .B(n204), .Y(N345));
sg13g2_nor2_2 U493 (.A(n184), .B(n204), .Y(N344));
sg13g2_inv_2 U494 (.A(n521), .Y(n1469));
sg13g2_inv_2 U495 (.A(n522), .Y(n1472));
sg13g2_inv_2 U496 (.A(n523), .Y(N462));
sg13g2_nand2_2 U497 (.A(n376), .B(n375), .Y(N341));
sg13g2_inv_2 U498 (.A(n524), .Y(n1477));
sg13g2_inv_2 U499 (.A(n525), .Y(n1478));
sg13g2_inv_2 U500 (.A(n526), .Y(n1481));
sg13g2_inv_2 U501 (.A(n527), .Y(N463));
sg13g2_nor2_2 U502 (.A(n391), .B(n392), .Y(n373));
sg13g2_nor2_2 U503 (.A(n379), .B(n204), .Y(N338));
sg13g2_inv_2 U504 (.A(n529), .Y(n1486));
sg13g2_nor2_2 U505 (.A(n204), .B(n380), .Y(N337));
sg13g2_nor2_2 U506 (.A(n380), .B(n376), .Y(N336));
sg13g2_inv_2 U507 (.A(n530), .Y(n1487));
sg13g2_inv_2 U508 (.A(n531), .Y(n1490));
sg13g2_inv_2 U509 (.A(n533), .Y(N464));
sg13g2_inv_2 U510 (.A(n535), .Y(n1495));
sg13g2_inv_2 U511 (.A(n536), .Y(n1496));
sg13g2_inv_2 U512 (.A(n537), .Y(n1499));
sg13g2_inv_2 U513 (.A(n539), .Y(N465));
sg13g2_inv_2 U514 (.A(n541), .Y(n1504));
sg13g2_inv_2 U515 (.A(n543), .Y(n1505));
sg13g2_inv_2 U516 (.A(n544), .Y(n1508));
sg13g2_inv_2 U517 (.A(n545), .Y(N466));
sg13g2_inv_2 U518 (.A(n546), .Y(n1513));
sg13g2_inv_2 U519 (.A(n547), .Y(n1514));
sg13g2_inv_2 U520 (.A(n548), .Y(n1517));
sg13g2_inv_2 U521 (.A(n552), .Y(N467));
sg13g2_inv_2 U522 (.A(n553), .Y(n1343));
sg13g2_inv_2 U523 (.A(n554), .Y(n1349));
sg13g2_inv_2 U524 (.A(n555), .Y(n1348));
sg13g2_inv_2 U525 (.A(n556), .Y(n1352));
sg13g2_inv_2 U526 (.A(n561), .Y(n1351));
sg13g2_inv_2 U527 (.A(n564), .Y(n1353));
sg13g2_inv_2 U528 (.A(n565), .Y(n1390));
sg13g2_inv_2 U529 (.A(n566), .Y(n1389));
sg13g2_inv_2 U530 (.A(n567), .Y(n1393));
sg13g2_nor2_2 U531 (.A(n372), .B(n128), .Y(N312));
sg13g2_nor2_2 U532 (.A(n372), .B(n132), .Y(N311));
sg13g2_nor2_2 U533 (.A(n372), .B(n136), .Y(N310));
sg13g2_nor2_2 U534 (.A(n372), .B(n140), .Y(N309));
sg13g2_nor2_2 U535 (.A(n372), .B(n144), .Y(N308));
sg13g2_nor2_2 U536 (.A(n372), .B(n148), .Y(N307));
sg13g2_nor2_2 U537 (.A(n372), .B(n152), .Y(N306));
sg13g2_nor2_2 U538 (.A(n372), .B(n156), .Y(N305));
sg13g2_nor2_2 U539 (.A(n372), .B(n184), .Y(N304));
sg13g2_inv_2 U540 (.A(n571), .Y(n1392));
sg13g2_inv_2 U541 (.A(n572), .Y(n1394));
sg13g2_nor2_2 U542 (.A(n207), .B(n381), .Y(N302));
sg13g2_inv_2 U543 (.A(n573), .Y(n1399));
sg13g2_nor2_2 U544 (.A(n211), .B(n381), .Y(N301));
sg13g2_inv_2 U545 (.A(n574), .Y(n1398));
sg13g2_nor2_2 U546 (.A(n213), .B(n381), .Y(N300));
sg13g2_inv_2 U547 (.A(n575), .Y(n1402));
sg13g2_nor2_2 U548 (.A(n215), .B(n381), .Y(N299));
sg13g2_inv_2 U549 (.A(n576), .Y(n1401));
sg13g2_nor2_2 U550 (.A(n217), .B(n381), .Y(N298));
sg13g2_inv_2 U551 (.A(n577), .Y(n1403));
sg13g2_nor2_2 U552 (.A(n219), .B(n381), .Y(N297));
sg13g2_inv_2 U553 (.A(n578), .Y(n1408));
sg13g2_nor2_2 U554 (.A(n221), .B(n381), .Y(N296));
sg13g2_inv_2 U555 (.A(n579), .Y(n1407));
sg13g2_nor2_2 U556 (.A(n223), .B(n381), .Y(N295));
sg13g2_inv_2 U557 (.A(n580), .Y(n1411));
sg13g2_nor2_2 U558 (.A(n225), .B(n381), .Y(N294));
sg13g2_inv_2 U559 (.A(n581), .Y(n1410));
sg13g2_nor2_2 U560 (.A(n227), .B(n381), .Y(N293));
sg13g2_inv_2 U561 (.A(n582), .Y(n1412));
sg13g2_inv_2 U562 (.A(n583), .Y(n1417));
sg13g2_inv_2 U563 (.A(n584), .Y(n1416));
sg13g2_nor2_2 U564 (.A(n231), .B(n381), .Y(N291));
sg13g2_inv_2 U565 (.A(n585), .Y(n1420));
sg13g2_nor2_2 U566 (.A(n233), .B(n381), .Y(N290));
sg13g2_inv_2 U567 (.A(n586), .Y(n1419));
sg13g2_nor2_2 U568 (.A(n235), .B(n381), .Y(N289));
sg13g2_inv_2 U569 (.A(n587), .Y(n1421));
sg13g2_nor2_2 U570 (.A(n237), .B(n381), .Y(N288));
sg13g2_inv_2 U571 (.A(n588), .Y(n1426));
sg13g2_nor2_2 U572 (.A(n239), .B(n381), .Y(N287));
sg13g2_inv_2 U573 (.A(n589), .Y(n1425));
sg13g2_nor2_2 U574 (.A(n160), .B(n381), .Y(N286));
sg13g2_inv_2 U575 (.A(n590), .Y(n1429));
sg13g2_nor2_2 U576 (.A(n164), .B(n381), .Y(N285));
sg13g2_inv_2 U577 (.A(n591), .Y(n1428));
sg13g2_nor2_2 U578 (.A(n168), .B(n381), .Y(N284));
sg13g2_inv_2 U579 (.A(n592), .Y(n1430));
sg13g2_nor2_2 U580 (.A(n172), .B(n381), .Y(N283));
sg13g2_inv_2 U581 (.A(n593), .Y(n1435));
sg13g2_nor2_2 U582 (.A(n176), .B(n381), .Y(N282));
sg13g2_inv_2 U583 (.A(n594), .Y(n1434));
sg13g2_nor2_2 U584 (.A(n180), .B(n381), .Y(N281));
sg13g2_inv_2 U585 (.A(n595), .Y(n1438));
sg13g2_nor2_2 U586 (.A(n124), .B(n381), .Y(N280));
sg13g2_inv_2 U587 (.A(n596), .Y(n1437));
sg13g2_nor2_2 U588 (.A(n128), .B(n381), .Y(N279));
sg13g2_inv_2 U589 (.A(n597), .Y(n1439));
sg13g2_nor2_2 U590 (.A(n132), .B(n381), .Y(N278));
sg13g2_inv_2 U591 (.A(sum_7), .Y(n132));
sg13g2_nor2_2 U592 (.A(n136), .B(n381), .Y(N277));
sg13g2_inv_2 U593 (.A(n598), .Y(n1444));
sg13g2_nor2_2 U594 (.A(n140), .B(n381), .Y(N276));
sg13g2_inv_2 U595 (.A(sum_5), .Y(n140));
sg13g2_nor2_2 U596 (.A(n144), .B(n381), .Y(N275));
sg13g2_inv_2 U597 (.A(sum_4), .Y(n144));
sg13g2_nor2_2 U598 (.A(n148), .B(n381), .Y(N274));
sg13g2_inv_2 U599 (.A(sum_3), .Y(n148));
sg13g2_nor2_2 U600 (.A(n152), .B(n381), .Y(N273));
sg13g2_inv_2 U601 (.A(sum_2), .Y(n152));
sg13g2_nor2_2 U602 (.A(n156), .B(n381), .Y(N272));
sg13g2_inv_2 U603 (.A(sum_1), .Y(n156));
sg13g2_nor2_2 U604 (.A(n184), .B(n381), .Y(N271));
sg13g2_inv_2 U605 (.A(sum_0), .Y(n184));
sg13g2_inv_2 U606 (.A(n599), .Y(n1443));
sg13g2_inv_2 U607 (.A(n600), .Y(n1447));
sg13g2_nand2_2 U608 (.A(n381), .B(n384), .Y(N269));
sg13g2_inv_2 U609 (.A(n385), .Y(N268));
sg13g2_inv_2 U610 (.A(n384), .Y(N259));
sg13g2_inv_2 U611 (.A(n601), .Y(n1446));
sg13g2_inv_2 U612 (.A(n602), .Y(n1448));
sg13g2_inv_2 U613 (.A(n603), .Y(n1453));
sg13g2_inv_2 U614 (.A(n604), .Y(n1452));
sg13g2_inv_2 U615 (.A(n605), .Y(n1456));
sg13g2_inv_2 U616 (.A(n606), .Y(n1455));
sg13g2_inv_2 U617 (.A(n607), .Y(n1457));
sg13g2_inv_2 U618 (.A(n608), .Y(n1462));
sg13g2_inv_2 U619 (.A(n609), .Y(n1461));
sg13g2_inv_2 U620 (.A(n610), .Y(n1465));
sg13g2_inv_2 U621 (.A(n611), .Y(n1464));
sg13g2_inv_2 U622 (.A(n399), .Y(n388));
sg13g2_inv_2 U623 (.A(n612), .Y(n1466));
sg13g2_inv_2 U624 (.A(n613), .Y(n1471));
sg13g2_inv_2 U625 (.A(n614), .Y(n1470));
sg13g2_inv_2 U626 (.A(n615), .Y(n1474));
sg13g2_nor2_2 U627 (.A(n392), .B(n393), .Y(n390));
sg13g2_inv_2 U628 (.A(n398), .Y(n389));
sg13g2_inv_2 U629 (.A(n616), .Y(n1473));
sg13g2_inv_2 U630 (.A(n617), .Y(n1475));
sg13g2_inv_2 U631 (.A(n618), .Y(n1558));
sg13g2_inv_2 U632 (.A(n619), .Y(n1480));
sg13g2_inv_2 U633 (.A(n620), .Y(n1479));
sg13g2_inv_2 U634 (.A(n621), .Y(n1483));
sg13g2_inv_2 U635 (.A(n622), .Y(n1482));
sg13g2_inv_2 U636 (.A(n623), .Y(n1484));
sg13g2_inv_2 U637 (.A(n624), .Y(n1559));
sg13g2_inv_2 U638 (.A(n625), .Y(n1489));
sg13g2_inv_2 U639 (.A(n626), .Y(n1488));
sg13g2_inv_2 U640 (.A(n627), .Y(n1492));
sg13g2_inv_2 U641 (.A(n628), .Y(n1491));
sg13g2_inv_2 U642 (.A(n629), .Y(n1493));
sg13g2_inv_2 U643 (.A(n630), .Y(n1560));
sg13g2_inv_2 U644 (.A(n631), .Y(n1498));
sg13g2_inv_2 U645 (.A(n632), .Y(n1497));
sg13g2_inv_2 U646 (.A(n633), .Y(n1501));
sg13g2_inv_2 U647 (.A(n634), .Y(n1500));
sg13g2_inv_2 U648 (.A(n635), .Y(n1502));
sg13g2_inv_2 U649 (.A(n636), .Y(n1561));
sg13g2_inv_2 U650 (.A(n637), .Y(n1507));
sg13g2_inv_2 U651 (.A(n638), .Y(n1506));
sg13g2_inv_2 U652 (.A(n639), .Y(n1510));
sg13g2_inv_2 U653 (.A(n640), .Y(n1509));
sg13g2_inv_2 U654 (.A(n641), .Y(n1511));
sg13g2_inv_2 U655 (.A(n642), .Y(n1562));
sg13g2_inv_2 U656 (.A(n643), .Y(n1516));
sg13g2_inv_2 U657 (.A(n644), .Y(n1515));
sg13g2_inv_2 U658 (.A(n645), .Y(n1519));
sg13g2_inv_2 U659 (.A(n646), .Y(n1518));
sg13g2_inv_2 U660 (.A(n647), .Y(n1520));
sg13g2_inv_2 U661 (.A(n648), .Y(n1563));
sg13g2_inv_2 U662 (.A(n649), .Y(n1566));
sg13g2_inv_2 U663 (.A(n650), .Y(n1564));
sg13g2_inv_2 U672 (.A(N135), .Y(n423));
sg13g2_inv_2 U678 (.A(N146), .Y(n429));
sg13g2_inv_2 U706 (.A(N200), .Y(n457));
sg13g2_inv_2 U801 (.A(n549), .Y(N541));
sg13g2_mux2_1 U822 (.A0(ki_0), .A1(\i_wb_data[0]), .S(N82), .X(n1103));
sg13g2_mux2_1 U824 (.A0(ki_1), .A1(\i_wb_data[1]), .S(N82), .X(n1102));
sg13g2_mux2_1 U826 (.A0(ki_2), .A1(\i_wb_data[2]), .S(N82), .X(n1101));
sg13g2_mux2_1 U828 (.A0(ki_3), .A1(\i_wb_data[3]), .S(N82), .X(n1100));
sg13g2_mux2_1 U830 (.A0(ki_4), .A1(\i_wb_data[4]), .S(N82), .X(n1099));
sg13g2_mux2_1 U832 (.A0(ki_5), .A1(\i_wb_data[5]), .S(N82), .X(n1098));
sg13g2_mux2_1 U834 (.A0(ki_6), .A1(\i_wb_data[6]), .S(N82), .X(n1097));
sg13g2_mux2_1 U836 (.A0(ki_7), .A1(\i_wb_data[7]), .S(N82), .X(n1096));
sg13g2_mux2_1 U838 (.A0(ki_8), .A1(\i_wb_data[8]), .S(N82), .X(n1095));
sg13g2_mux2_1 U840 (.A0(ki_9), .A1(\i_wb_data[9]), .S(N82), .X(n1094));
sg13g2_mux2_1 U842 (.A0(ki_10), .A1(\i_wb_data[10]), .S(N82), .X(n1093));
sg13g2_mux2_1 U844 (.A0(ki_11), .A1(\i_wb_data[11]), .S(N82), .X(n1092));
sg13g2_mux2_1 U846 (.A0(ki_12), .A1(\i_wb_data[12]), .S(N82), .X(n1091));
sg13g2_mux2_1 U848 (.A0(ki_13), .A1(\i_wb_data[13]), .S(N82), .X(n1090));
sg13g2_mux2_1 U850 (.A0(ki_14), .A1(\i_wb_data[14]), .S(N82), .X(n1089));
sg13g2_mux2_1 U852 (.A0(ki_15), .A1(\i_wb_data[15]), .S(N82), .X(n1088));
sg13g2_mux2_1 U854 (.A0(kd_0), .A1(\i_wb_data[0]), .S(N85), .X(n1087));
sg13g2_mux2_1 U856 (.A0(kd_1), .A1(\i_wb_data[1]), .S(N85), .X(n1086));
sg13g2_mux2_1 U858 (.A0(kd_2), .A1(\i_wb_data[2]), .S(N85), .X(n1085));
sg13g2_mux2_1 U860 (.A0(kd_3), .A1(\i_wb_data[3]), .S(N85), .X(n1084));
sg13g2_mux2_1 U862 (.A0(kd_4), .A1(\i_wb_data[4]), .S(N85), .X(n1083));
sg13g2_mux2_1 U864 (.A0(kd_5), .A1(\i_wb_data[5]), .S(N85), .X(n1082));
sg13g2_mux2_1 U866 (.A0(kd_6), .A1(\i_wb_data[6]), .S(N85), .X(n1081));
sg13g2_mux2_1 U868 (.A0(kd_7), .A1(\i_wb_data[7]), .S(N85), .X(n1080));
sg13g2_mux2_1 U870 (.A0(kd_8), .A1(\i_wb_data[8]), .S(N85), .X(n1079));
sg13g2_mux2_1 U872 (.A0(kd_9), .A1(\i_wb_data[9]), .S(N85), .X(n1078));
sg13g2_mux2_1 U874 (.A0(kd_10), .A1(\i_wb_data[10]), .S(N85), .X(n1077));
sg13g2_mux2_1 U876 (.A0(kd_11), .A1(\i_wb_data[11]), .S(N85), .X(n1076));
sg13g2_mux2_1 U878 (.A0(kd_12), .A1(\i_wb_data[12]), .S(N85), .X(n1075));
sg13g2_mux2_1 U880 (.A0(kd_13), .A1(\i_wb_data[13]), .S(N85), .X(n1074));
sg13g2_mux2_1 U882 (.A0(kd_14), .A1(\i_wb_data[14]), .S(N85), .X(n1073));
sg13g2_mux2_1 U884 (.A0(kd_15), .A1(\i_wb_data[15]), .S(N85), .X(n1072));
sg13g2_mux2_1 U886 (.A0(sp_0), .A1(\i_wb_data[0]), .S(N86), .X(n1071));
sg13g2_mux2_1 U888 (.A0(sp_1), .A1(\i_wb_data[1]), .S(N86), .X(n1070));
sg13g2_mux2_1 U890 (.A0(sp_2), .A1(\i_wb_data[2]), .S(N86), .X(n1069));
sg13g2_mux2_1 U892 (.A0(sp_3), .A1(\i_wb_data[3]), .S(N86), .X(n1068));
sg13g2_mux2_1 U894 (.A0(sp_4), .A1(\i_wb_data[4]), .S(N86), .X(n1067));
sg13g2_mux2_1 U896 (.A0(sp_5), .A1(\i_wb_data[5]), .S(N86), .X(n1066));
sg13g2_mux2_1 U898 (.A0(sp_6), .A1(\i_wb_data[6]), .S(N86), .X(n1065));
sg13g2_mux2_1 U900 (.A0(sp_7), .A1(\i_wb_data[7]), .S(N86), .X(n1064));
sg13g2_mux2_1 U902 (.A0(sp_8), .A1(\i_wb_data[8]), .S(N86), .X(n1063));
sg13g2_mux2_1 U904 (.A0(sp_9), .A1(\i_wb_data[9]), .S(N86), .X(n1062));
sg13g2_mux2_1 U906 (.A0(sp_10), .A1(\i_wb_data[10]), .S(N86), .X(n1061));
sg13g2_mux2_1 U908 (.A0(sp_11), .A1(\i_wb_data[11]), .S(N86), .X(n1060));
sg13g2_mux2_1 U910 (.A0(sp_12), .A1(\i_wb_data[12]), .S(N86), .X(n1059));
sg13g2_mux2_1 U912 (.A0(sp_13), .A1(\i_wb_data[13]), .S(N86), .X(n1058));
sg13g2_mux2_1 U914 (.A0(sp_14), .A1(\i_wb_data[14]), .S(N86), .X(n1057));
sg13g2_mux2_1 U916 (.A0(sp_15), .A1(\i_wb_data[15]), .S(N86), .X(n1056));
sg13g2_mux2_1 U918 (.A0(pv_0), .A1(\i_wb_data[0]), .S(N87), .X(n1055));
sg13g2_mux2_1 U920 (.A0(pv_1), .A1(\i_wb_data[1]), .S(N87), .X(n1054));
sg13g2_mux2_1 U922 (.A0(pv_2), .A1(\i_wb_data[2]), .S(N87), .X(n1053));
sg13g2_mux2_1 U924 (.A0(pv_3), .A1(\i_wb_data[3]), .S(N87), .X(n1052));
sg13g2_mux2_1 U926 (.A0(pv_4), .A1(\i_wb_data[4]), .S(N87), .X(n1051));
sg13g2_mux2_1 U928 (.A0(pv_5), .A1(\i_wb_data[5]), .S(N87), .X(n1050));
sg13g2_mux2_1 U930 (.A0(pv_6), .A1(\i_wb_data[6]), .S(N87), .X(n1049));
sg13g2_mux2_1 U932 (.A0(pv_7), .A1(\i_wb_data[7]), .S(N87), .X(n1048));
sg13g2_mux2_1 U934 (.A0(pv_8), .A1(\i_wb_data[8]), .S(N87), .X(n1047));
sg13g2_mux2_1 U936 (.A0(pv_9), .A1(\i_wb_data[9]), .S(N87), .X(n1046));
sg13g2_mux2_1 U938 (.A0(pv_10), .A1(\i_wb_data[10]), .S(N87), .X(n1045));
sg13g2_mux2_1 U940 (.A0(pv_11), .A1(\i_wb_data[11]), .S(N87), .X(n1044));
sg13g2_mux2_1 U942 (.A0(pv_12), .A1(\i_wb_data[12]), .S(N87), .X(n1043));
sg13g2_mux2_1 U944 (.A0(pv_13), .A1(\i_wb_data[13]), .S(N87), .X(n1042));
sg13g2_mux2_1 U946 (.A0(pv_14), .A1(\i_wb_data[14]), .S(N87), .X(n1041));
sg13g2_mux2_1 U948 (.A0(pv_15), .A1(\i_wb_data[15]), .S(N87), .X(n1040));
sg13g2_mux2_1 U950 (.A0(kp_0), .A1(\i_wb_data[0]), .S(N88), .X(n1039));
sg13g2_mux2_1 U952 (.A0(kp_1), .A1(\i_wb_data[1]), .S(N88), .X(n1038));
sg13g2_mux2_1 U954 (.A0(kp_2), .A1(\i_wb_data[2]), .S(N88), .X(n1037));
sg13g2_mux2_1 U956 (.A0(kp_3), .A1(\i_wb_data[3]), .S(N88), .X(n1036));
sg13g2_mux2_1 U958 (.A0(kp_4), .A1(\i_wb_data[4]), .S(N88), .X(n1035));
sg13g2_mux2_1 U960 (.A0(kp_5), .A1(\i_wb_data[5]), .S(N88), .X(n1034));
sg13g2_mux2_1 U962 (.A0(kp_6), .A1(\i_wb_data[6]), .S(N88), .X(n1033));
sg13g2_mux2_1 U964 (.A0(kp_7), .A1(\i_wb_data[7]), .S(N88), .X(n1032));
sg13g2_mux2_1 U966 (.A0(kp_8), .A1(\i_wb_data[8]), .S(N88), .X(n1031));
sg13g2_mux2_1 U968 (.A0(kp_9), .A1(\i_wb_data[9]), .S(N88), .X(n1030));
sg13g2_mux2_1 U970 (.A0(kp_10), .A1(\i_wb_data[10]), .S(N88), .X(n1029));
sg13g2_mux2_1 U972 (.A0(kp_11), .A1(\i_wb_data[11]), .S(N88), .X(n1028));
sg13g2_mux2_1 U974 (.A0(kp_12), .A1(\i_wb_data[12]), .S(N88), .X(n1027));
sg13g2_mux2_1 U976 (.A0(kp_13), .A1(\i_wb_data[13]), .S(N88), .X(n1026));
sg13g2_mux2_1 U978 (.A0(kp_14), .A1(\i_wb_data[14]), .S(N88), .X(n1025));
sg13g2_mux2_1 U980 (.A0(kp_15), .A1(\i_wb_data[15]), .S(N88), .X(n1024));
sg13g2_mux2_1 U1002 (.A0(cout), .A1(n396), .S(N426), .X(n1013));
sg13g2_mux2_1 U1004 (.A0(start), .A1(n396), .S(N427), .X(n1012));
sg13g2_mux2_1 U1006 (.A0(rl_5), .A1(n399), .S(N268), .X(n1011));
sg13g2_mux2_1 U1020 (.A0(p_0), .A1(N361), .S(net9475), .X(n1004));
sg13g2_mux2_1 U1022 (.A0(p_1), .A1(N362), .S(net9476), .X(n1003));
sg13g2_mux2_1 U1024 (.A0(p_2), .A1(N363), .S(net9475), .X(n1002));
sg13g2_mux2_1 U1026 (.A0(p_3), .A1(N364), .S(net9476), .X(n1001));
sg13g2_mux2_1 U1028 (.A0(p_4), .A1(N365), .S(net9475), .X(n1000));
sg13g2_mux2_1 U1030 (.A0(p_5), .A1(N366), .S(net9476), .X(n999));
sg13g2_mux2_1 U1032 (.A0(p_6), .A1(N367), .S(net9475), .X(n998));
sg13g2_mux2_1 U1034 (.A0(p_7), .A1(N368), .S(net9476), .X(n997));
sg13g2_mux2_1 U1036 (.A0(p_8), .A1(N369), .S(net9475), .X(n996));
sg13g2_mux2_1 U1038 (.A0(p_9), .A1(N370), .S(net9476), .X(n995));
sg13g2_mux2_1 U1040 (.A0(p_10), .A1(N371), .S(net9475), .X(n994));
sg13g2_mux2_1 U1042 (.A0(p_11), .A1(N372), .S(net9476), .X(n993));
sg13g2_mux2_1 U1046 (.A0(p_13), .A1(N374), .S(net9476), .X(n991));
sg13g2_mux2_1 U1050 (.A0(p_15), .A1(N376), .S(net9476), .X(n989));
sg13g2_mux2_1 U1062 (.A0(p_21), .A1(n1310), .S(net9476), .X(n983));
sg13g2_mux2_1 U1148 (.A0(\o_un[0]), .A1(N271), .S(N270), .X(n940));
sg13g2_mux2_1 U1150 (.A0(\o_un[1]), .A1(N272), .S(N270), .X(n939));
sg13g2_mux2_1 U1152 (.A0(\o_un[2]), .A1(N273), .S(N270), .X(n938));
sg13g2_mux2_1 U1154 (.A0(\o_un[3]), .A1(N274), .S(N270), .X(n937));
sg13g2_mux2_1 U1156 (.A0(\o_un[4]), .A1(N275), .S(N270), .X(n936));
sg13g2_mux2_1 U1158 (.A0(\o_un[5]), .A1(N276), .S(N270), .X(n935));
sg13g2_mux2_1 U1160 (.A0(\o_un[6]), .A1(N277), .S(N270), .X(n934));
sg13g2_mux2_1 U1162 (.A0(\o_un[7]), .A1(N278), .S(N270), .X(n933));
sg13g2_mux2_1 U1164 (.A0(\o_un[8]), .A1(N279), .S(N270), .X(n932));
sg13g2_mux2_1 U1166 (.A0(\o_un[9]), .A1(N280), .S(N270), .X(n931));
sg13g2_mux2_1 U1168 (.A0(\o_un[10]), .A1(N281), .S(N270), .X(n930));
sg13g2_mux2_1 U1170 (.A0(\o_un[11]), .A1(N282), .S(N270), .X(n929));
sg13g2_mux2_1 U1172 (.A0(\o_un[12]), .A1(N283), .S(N270), .X(n928));
sg13g2_mux2_1 U1174 (.A0(\o_un[13]), .A1(N284), .S(N270), .X(n927));
sg13g2_mux2_1 U1176 (.A0(\o_un[14]), .A1(N285), .S(N270), .X(n926));
sg13g2_mux2_1 U1178 (.A0(\o_un[15]), .A1(N286), .S(N270), .X(n925));
sg13g2_mux2_1 U1180 (.A0(\o_un[16]), .A1(N287), .S(N270), .X(n924));
sg13g2_mux2_1 U1182 (.A0(\o_un[17]), .A1(N288), .S(N270), .X(n923));
sg13g2_mux2_1 U1184 (.A0(\o_un[18]), .A1(N289), .S(N270), .X(n922));
sg13g2_mux2_1 U1186 (.A0(\o_un[19]), .A1(N290), .S(N270), .X(n921));
sg13g2_mux2_1 U1188 (.A0(\o_un[20]), .A1(N291), .S(N270), .X(n920));
sg13g2_mux2_1 U1190 (.A0(\o_un[21]), .A1(N292), .S(N270), .X(n919));
sg13g2_mux2_1 U1194 (.A0(\o_un[23]), .A1(N294), .S(N270), .X(n917));
sg13g2_mux2_1 U1196 (.A0(\o_un[24]), .A1(N295), .S(N270), .X(n916));
sg13g2_mux2_1 U1198 (.A0(\o_un[25]), .A1(N296), .S(N270), .X(n915));
sg13g2_mux2_1 U1200 (.A0(\o_un[26]), .A1(N297), .S(N270), .X(n914));
sg13g2_mux2_1 U1202 (.A0(\o_un[27]), .A1(N298), .S(N270), .X(n913));
sg13g2_mux2_1 U1204 (.A0(\o_un[28]), .A1(N299), .S(N270), .X(n912));
sg13g2_mux2_1 U1206 (.A0(\o_un[29]), .A1(N300), .S(N270), .X(n911));
sg13g2_mux2_1 U1208 (.A0(\o_un[30]), .A1(N301), .S(N270), .X(n910));
sg13g2_mux2_1 U1210 (.A0(\o_un[31]), .A1(N302), .S(N270), .X(n909));
sg13g2_mux2_1 U1222 (.A0(sigma_5), .A1(N309), .S(n1313), .X(n903));
sg13g2_mux2_1 U1224 (.A0(sigma_6), .A1(N310), .S(n1313), .X(n902));
sg13g2_mux2_1 U1226 (.A0(sigma_7), .A1(N311), .S(n1313), .X(n901));
sg13g2_mux2_1 U1230 (.A0(sigma_9), .A1(N313), .S(n1313), .X(n899));
sg13g2_mux2_1 U1232 (.A0(sigma_10), .A1(N314), .S(n1313), .X(n898));
sg13g2_mux2_1 U1234 (.A0(sigma_11), .A1(N315), .S(n1313), .X(n897));
sg13g2_mux2_1 U1238 (.A0(sigma_13), .A1(N317), .S(n1313), .X(n895));
sg13g2_mux2_1 U1244 (.A0(sigma_16), .A1(N320), .S(n1313), .X(n892));
sg13g2_mux2_1 U1246 (.A0(sigma_17), .A1(N321), .S(n1313), .X(n891));
sg13g2_mux2_1 U1250 (.A0(sigma_19), .A1(N323), .S(n1313), .X(n889));
sg13g2_mux2_1 U1254 (.A0(sigma_21), .A1(N325), .S(n1313), .X(n887));
sg13g2_mux2_1 U1270 (.A0(sigma_29), .A1(N333), .S(n1313), .X(n879));
sg13g2_mux2_1 U1274 (.A0(sigma_31), .A1(N335), .S(n1313), .X(n877));
sg13g2_mux2_1 U1276 (.A0(a_0), .A1(N393), .S(net9475), .X(n876));
sg13g2_mux2_1 U1278 (.A0(a_1), .A1(N394), .S(net9476), .X(n875));
sg13g2_mux2_1 U1280 (.A0(a_2), .A1(N395), .S(net9475), .X(n874));
sg13g2_mux2_1 U1282 (.A0(a_3), .A1(N396), .S(net9476), .X(n873));
sg13g2_mux2_1 U1284 (.A0(a_4), .A1(N397), .S(net9475), .X(n872));
sg13g2_mux2_1 U1286 (.A0(a_5), .A1(N398), .S(net9476), .X(n871));
sg13g2_mux2_1 U1288 (.A0(a_6), .A1(N399), .S(net9475), .X(n870));
sg13g2_mux2_1 U1290 (.A0(a_7), .A1(N400), .S(net9476), .X(n869));
sg13g2_mux2_1 U1294 (.A0(a_9), .A1(N402), .S(net9476), .X(n867));
sg13g2_mux2_1 U1296 (.A0(a_10), .A1(N403), .S(net9475), .X(n866));
sg13g2_mux2_1 U1298 (.A0(a_11), .A1(N404), .S(net9476), .X(n865));
sg13g2_mux2_1 U1312 (.A0(of_0), .A1(N336), .S(N341), .X(n858));
sg13g2_mux2_1 U1316 (.A0(a_17), .A1(N410), .S(net9476), .X(n856));
sg13g2_nor2_2 U1484 (.A(n211), .B(n372), .Y(n1241));
sg13g2_mux2_1 U1485 (.A0(\o_un[22]), .A1(N293), .S(N270), .X(n918));
sg13g2_nand3_1 U1487 (.A(n320), .B(n321), .C(n322), .Y(N373));
sg13g2_nand2_2 U1488 (.A(product_12), .B(n292), .Y(n321));
sg13g2_a21oi_2 U1490 (.A1(sigma_27), .A2(N263), .B1(N331), .Y(n218));
sg13g2_o21ai_1 U1491 (.A1(of_4), .A2(\of_addition[1]), .B1(n393), .Y(n377));
sg13g2_mux2_1 U1492 (.A0(N424), .A1(a_31), .S(n1242), .X(n842));
sg13g2_inv_2 U1493 (.A(net9476), .Y(n1242));
sg13g2_mux2_1 U1494 (.A0(a_19), .A1(N412), .S(net9476), .X(n854));
sg13g2_mux2_1 U1495 (.A0(N379), .A1(p_18), .S(net14608), .X(n986));
sg13g2_nand2_2 U1496 (.A(product_14), .B(n292), .Y(n313));
sg13g2_mux2_1 U1497 (.A0(p_14), .A1(N375), .S(net9475), .X(n990));
sg13g2_mux2_1 U1498 (.A0(sigma_14), .A1(N318), .S(n1313), .X(n894));
sg13g2_a21oi_2 U1499 (.A1(n398), .A2(kd_14), .B1(N318), .Y(n244));
sg13g2_nor2_2 U1500 (.A(n372), .B(n164), .Y(N318));
sg13g2_mux2_1 U1501 (.A0(n1308), .A1(p_27), .S(n1297), .X(n977));
sg13g2_mux2_1 U1502 (.A0(net9913), .A1(n294), .S(net9475), .X(n443));
sg13g2_a21oi_2 U1503 (.A1(product_29), .A2(n292), .B1(n293), .Y(n295));
sg13g2_a21oi_2 U1504 (.A1(product_20), .A2(n292), .B1(n293), .Y(n304));
sg13g2_mux2_1 U1505 (.A0(n1304), .A1(n304), .S(N360), .X(n447));
sg13g2_o21ai_1 U1506 (.A1(pv_15), .A2(n206), .B1(n243), .Y(n242));
sg13g2_inv_2 U1507 (.A(net9474), .Y(net9475));
sg13g2_inv_2 U1508 (.A(n1321), .Y(n1322));
sg13g2_inv_2 U1509 (.A(N190), .Y(n452));
sg13g2_a21oi_2 U1512 (.A1(sigma_23), .A2(N263), .B1(N327), .Y(n226));
sg13g2_inv_2 U1514 (.A(N303), .Y(n374));
sg13g2_inv_2 U1515 (.A(net14330), .Y(n1296));
sg13g2_a21oi_2 U1518 (.A1(sigma_28), .A2(N263), .B1(N332), .Y(n216));
sg13g2_a21oi_2 U1520 (.A1(sigma_31), .A2(N263), .B1(N335), .Y(n210));
sg13g2_inv_2 U1530 (.A(net9476), .Y(net13458));
sg13g2_inv_2 U1538 (.A(net9476), .Y(n1297));
sg13g2_nand2_2 U1575 (.A(state_1_4), .B(N150), .Y(n1243));
sg13g2_inv_2 U1576 (.A(n1243), .Y(n426));
sg13g2_nor2_2 U1578 (.A(N151), .B(N174), .Y(n444));
sg13g2_nand3_1 U1579 (.A(n190), .B(n199), .C(n1525), .Y(n1244));
sg13g2_inv_2 U1580 (.A(n1244), .Y(N87));
sg13g2_mux2_1 U1581 (.A0(sigma_4), .A1(N308), .S(n1313), .X(n904));
sg13g2_nand2_2 U1583 (.A(N139), .B(state_1_5), .Y(N153));
sg13g2_nand3_1 U1584 (.A(n446), .B(N183), .C(n431), .Y(N112));
sg13g2_nand2_2 U1587 (.A(N106), .B(N95), .Y(N177));
sg13g2_a21oi_2 U1588 (.A1(n1246), .A2(sigma_14), .B1(n246), .Y(n245));
sg13g2_inv_2 U1589 (.A(n1314), .Y(n1246));
sg13g2_mux2_1 U1590 (.A0(\err[0][4]), .A1(N348), .S(N342), .X(n952));
sg13g2_nor2_2 U1592 (.A(n1248), .B(md_index_1), .Y(N473));
sg13g2_nand2_2 U1594 (.A(N128), .B(N117), .Y(N198));
sg13g2_nor2_2 U1596 (.A(n388), .B(n36), .Y(N257));
sg13g2_nor2_2 U1597 (.A(n1318), .B(state_1_0), .Y(n1319));
sg13g2_mux2_1 U1599 (.A0(sigma_3), .A1(N307), .S(n1313), .X(n905));
sg13g2_nand3_1 U1601 (.A(n1525), .B(N480), .C(\i_wb_adr[4]), .Y(N520));
sg13g2_nand2_2 U1602 (.A(n402), .B(n456), .Y(N179));
sg13g2_inv_2 U1603 (.A(N98), .Y(n402));
sg13g2_nor2_2 U1604 (.A(state_1_7), .B(state_1_5), .Y(n1320));
sg13g2_mux2_1 U1606 (.A0(\err[0][3]), .A1(N347), .S(N342), .X(n953));
sg13g2_nor2_2 U1608 (.A(n1251), .B(md_index_0), .Y(N470));
sg13g2_nand2_2 U1610 (.A(n430), .B(n413), .Y(n1252));
sg13g2_inv_2 U1611 (.A(n1252), .Y(n416));
sg13g2_nand4_1 U1612 (.A(n399), .B(n36), .C(N542), .D(adr_check), .Y(n384));
sg13g2_nand4_1 U1613 (.A(N95), .B(n410), .C(n445), .D(state_1_1), .Y(n1262));
sg13g2_inv_2 U1614 (.A(N112), .Y(n410));
sg13g2_inv_2 U1615 (.A(N179), .Y(n445));
sg13g2_nand4_1 U1616 (.A(n1525), .B(n1341), .C(N480), .D(n190), .Y(n1253));
sg13g2_inv_2 U1617 (.A(n1253), .Y(N88));
sg13g2_mux2_1 U1619 (.A0(sigma_2), .A1(N306), .S(n1313), .X(n906));
sg13g2_nor2_2 U1621 (.A(state_1_8), .B(state_1_9), .Y(n1255));
sg13g2_inv_2 U1622 (.A(n1255), .Y(n1318));
sg13g2_nand2_2 U1623 (.A(n426), .B(n456), .Y(N146));
sg13g2_o21ai_1 U1624 (.A1(n1342), .A2(n1343), .B1(n1256), .Y(n568));
sg13g2_inv_2 U1625 (.A(n569), .Y(n1256));
sg13g2_nand3_1 U1626 (.A(n416), .B(n402), .C(n415), .Y(N125));
sg13g2_nor2_2 U1627 (.A(wlRS), .B(N484), .Y(N539));
sg13g2_nand3_1 U1628 (.A(n190), .B(n1525), .C(n200), .Y(n1257));
sg13g2_inv_2 U1629 (.A(n1257), .Y(N85));
sg13g2_mux2_1 U1630 (.A0(state_1_3), .A1(N259), .S(N255), .X(n1019));
sg13g2_mux2_1 U1633 (.A0(\err[0][2]), .A1(N346), .S(N342), .X(n954));
sg13g2_nor2_2 U1635 (.A(n1260), .B(\i_wb_data[8]), .Y(n508));
sg13g2_inv_2 U1636 (.A(n1336), .Y(n1260));
sg13g2_nand2_2 U1637 (.A(N172), .B(N161), .Y(n1261));
sg13g2_inv_2 U1638 (.A(n1261), .Y(n413));
sg13g2_nor2_2 U1641 (.A(md_index_1), .B(md_index_0), .Y(n1272));
sg13g2_inv_2 U1642 (.A(n1262), .Y(n398));
sg13g2_nand2_2 U1643 (.A(n430), .B(n431), .Y(N156));
sg13g2_nor2_2 U1644 (.A(\i_wb_adr[4]), .B(\i_wb_adr[3]), .Y(n1274));
sg13g2_nand4_1 U1645 (.A(N537), .B(i_wb_cyc), .C(i_wb_we), .D(i_wb_stb), .Y(n38));
sg13g2_mux2_1 U1647 (.A0(sigma_1), .A1(N305), .S(N303), .X(n907));
sg13g2_mux2_1 U1649 (.A0(\wl[0]), .A1(n399), .S(N266), .X(n1106));
sg13g2_nand3_1 U1651 (.A(n465), .B(n463), .C(n1329), .Y(N488));
sg13g2_nor2_2 U1652 (.A(\i_wb_data[22]), .B(n1288), .Y(n1265));
sg13g2_inv_2 U1653 (.A(n1265), .Y(N494));
sg13g2_nand3_1 U1654 (.A(n1266), .B(n493), .C(n1333), .Y(N503));
sg13g2_inv_2 U1655 (.A(\i_wb_data[13]), .Y(n1266));
sg13g2_nand3_1 U1656 (.A(n528), .B(n1335), .C(n1267), .Y(N525));
sg13g2_inv_2 U1657 (.A(\i_wb_adr[13]), .Y(n1267));
sg13g2_a21oi_2 U1658 (.A1(rl_6), .A2(\i_wb_adr[5]), .B1(rl_5), .Y(n1522));
sg13g2_nand2_2 U1659 (.A(p_31), .B(a_31), .Y(n1268));
sg13g2_inv_2 U1660 (.A(n1268), .Y(N554));
sg13g2_nand3_1 U1661 (.A(state_1_8), .B(n446), .C(n413), .Y(n1269));
sg13g2_inv_2 U1662 (.A(n1269), .Y(n451));
sg13g2_nand4_1 U1663 (.A(n508), .B(n511), .C(n1270), .D(n507), .Y(n1271));
sg13g2_inv_2 U1664 (.A(\i_wb_data[6]), .Y(n1270));
sg13g2_inv_2 U1665 (.A(n1271), .Y(n514));
sg13g2_nor2_2 U1666 (.A(state_1_7), .B(state_1_6), .Y(n431));
sg13g2_a21oi_2 U1667 (.A1(md_index_1), .A2(md_index_0), .B1(n1272), .Y(n123));
sg13g2_a21oi_2 U1668 (.A1(N547), .A2(n160), .B1(n1273), .Y(n380));
sg13g2_inv_2 U1669 (.A(n558), .Y(n1273));
sg13g2_nand2_2 U1670 (.A(N106), .B(N95), .Y(N122));
sg13g2_nand3_1 U1672 (.A(\i_wb_adr[2]), .B(n190), .C(n1274), .Y(n1275));
sg13g2_inv_2 U1673 (.A(n1275), .Y(N82));
sg13g2_inv_2 U1675 (.A(i_wb_stb), .Y(n1276));
sg13g2_mux2_1 U1676 (.A0(state_1_5), .A1(n395), .S(N255), .X(n1017));
sg13g2_nand4_1 U1679 (.A(state_0), .B(n1339), .C(n40), .D(N539), .Y(n1278));
sg13g2_inv_2 U1680 (.A(n1278), .Y(N81));
sg13g2_mux2_1 U1681 (.A0(wl_3), .A1(n399), .S(N269), .X(n1010));
sg13g2_nor2_2 U1683 (.A(n1280), .B(\i_wb_data[26]), .Y(n472));
sg13g2_inv_2 U1684 (.A(n1330), .Y(n1280));
sg13g2_nand3_1 U1685 (.A(n483), .B(n481), .C(n1331), .Y(N497));
sg13g2_nand3_1 U1686 (.A(n534), .B(n532), .C(n1337), .Y(N528));
sg13g2_nand4_1 U1687 (.A(N183), .B(N172), .C(N161), .D(state_1_9), .Y(N200));
sg13g2_nand3_1 U1688 (.A(i_wb_cyc), .B(i_wb_stb), .C(N534), .Y(n1281));
sg13g2_inv_2 U1689 (.A(n1281), .Y(re));
sg13g2_nor2_2 U1690 (.A(n1282), .B(mr_index_1), .Y(N476));
sg13g2_inv_2 U1691 (.A(mr_index_0), .Y(n1282));
sg13g2_nand4_1 U1692 (.A(n1341), .B(\i_wb_adr[2]), .C(\i_wb_adr[3]), .D(\i_wb_adr[5]), .Y(N484));
sg13g2_nor2_2 U1693 (.A(of_3), .B(\of_addition[1]), .Y(n378));
sg13g2_nand2_2 U1694 (.A(n432), .B(n456), .Y(N157));
sg13g2_nor2_2 U1695 (.A(\i_wb_data[1]), .B(N514), .Y(n1283));
sg13g2_inv_2 U1696 (.A(n1283), .Y(N515));
sg13g2_nand3_1 U1697 (.A(\i_wb_adr[2]), .B(n190), .C(n200), .Y(n1284));
sg13g2_inv_2 U1698 (.A(n1284), .Y(N86));
sg13g2_o21ai_1 U1699 (.A1(n123), .A2(n172), .B1(n173), .Y(md_12));
sg13g2_a21oi_2 U1700 (.A1(n1285), .A2(sigma_26), .B1(N330), .Y(n220));
sg13g2_inv_2 U1701 (.A(n1314), .Y(n1285));
sg13g2_nand3_1 U1702 (.A(n316), .B(n317), .C(n318), .Y(N374));
sg13g2_nand3_1 U1703 (.A(n324), .B(n325), .C(n326), .Y(N372));
sg13g2_nand3_1 U1704 (.A(n332), .B(n333), .C(n334), .Y(N370));
sg13g2_nand3_1 U1705 (.A(n336), .B(n337), .C(n338), .Y(N369));
sg13g2_nand3_1 U1706 (.A(n344), .B(n345), .C(n346), .Y(N367));
sg13g2_nand3_1 U1707 (.A(n352), .B(n353), .C(n354), .Y(N365));
sg13g2_mux2_1 U1709 (.A0(\err[0][1]), .A1(N345), .S(N342), .X(n955));
sg13g2_mux2_1 U1711 (.A0(rl_6), .A1(n399), .S(N269), .X(n1009));
sg13g2_o21ai_1 U1712 (.A1(N537), .A2(N536), .B1(n194), .Y(n1105));
sg13g2_nand4_1 U1713 (.A(n472), .B(n475), .C(n1287), .D(n471), .Y(n1288));
sg13g2_inv_2 U1714 (.A(\i_wb_data[24]), .Y(n1287));
sg13g2_nand3_1 U1715 (.A(n489), .B(n487), .C(n1332), .Y(N500));
sg13g2_nand3_1 U1716 (.A(n501), .B(n499), .C(n1334), .Y(N506));
sg13g2_nand2_2 U1717 (.A(N150), .B(N139), .Y(N98));
sg13g2_nand3_1 U1718 (.A(n540), .B(n538), .C(n1338), .Y(N531));
sg13g2_xnor2_1 U1719 (.A(mr_index_1), .B(mr_index_0), .Y(N91));
sg13g2_nor2_2 U1720 (.A(\wl[0]), .B(wl_3), .Y(n1289));
sg13g2_inv_2 U1721 (.A(n1289), .Y(wlRS));
sg13g2_nand4_1 U1722 (.A(n517), .B(n1290), .C(n513), .D(n514), .Y(N514));
sg13g2_inv_2 U1723 (.A(\i_wb_data[3]), .Y(n1290));
sg13g2_nor2_2 U1724 (.A(\i_wb_adr[3]), .B(\i_wb_adr[4]), .Y(n1530));
sg13g2_nor2_2 U1725 (.A(N188), .B(N191), .Y(n1291));
sg13g2_inv_2 U1726 (.A(n1291), .Y(n208));
sg13g2_inv_2 U1727 (.A(N153), .Y(n432));
sg13g2_o21ai_1 U1728 (.A1(n123), .A2(n160), .B1(n161), .Y(md_15));
sg13g2_a21oi_2 U1729 (.A1(n1292), .A2(sigma_18), .B1(N322), .Y(n236));
sg13g2_inv_2 U1730 (.A(n1314), .Y(n1292));
sg13g2_nand3_1 U1731 (.A(n340), .B(n341), .C(n342), .Y(N368));
sg13g2_nand3_1 U1732 (.A(n348), .B(n349), .C(n350), .Y(N366));
sg13g2_nand3_1 U1733 (.A(n356), .B(n357), .C(n358), .Y(N364));
sg13g2_nand3_1 U1734 (.A(n360), .B(n361), .C(n362), .Y(N363));
sg13g2_nand3_1 U1735 (.A(n364), .B(n365), .C(n366), .Y(N362));
sg13g2_mux2_1 U1736 (.A0(sigma_0), .A1(N304), .S(N303), .X(n908));
sg13g2_nand3_1 U1738 (.A(n368), .B(n369), .C(n370), .Y(N361));
sg13g2_xnor2_1 U1740 (.A(state_0), .B(N79), .Y(n1295));
sg13g2_inv_2 U1741 (.A(n1295), .Y(n1104));
sg13g2_inv_2 U1742 (.A(N151), .Y(n430));
sg13g2_inv_2 U1743 (.A(n1314), .Y(N263));
sg13g2_nand4_1 U1744 (.A(n1324), .B(n1323), .C(n1320), .D(n1319), .Y(n1314));
sg13g2_nand2_2 U1745 (.A(n381), .B(n375), .Y(N270));
sg13g2_nor2_2 U1746 (.A(N188), .B(N191), .Y(n392));
sg13g2_inv_2 U1747 (.A(n1), .Y(N430));
sg13g2_inv_2 U1748 (.A(N198), .Y(n456));
sg13g2_nor2_2 U1749 (.A(N100), .B(N103), .Y(n399));
sg13g2_inv_2 U1750 (.A(sum_15), .Y(n160));
sg13g2_nor2_2 U1752 (.A(N177), .B(N180), .Y(n393));
sg13g2_nor2_2 U1753 (.A(N122), .B(N125), .Y(n397));
sg13g2_nor2_2 U1754 (.A(N133), .B(N136), .Y(n396));
sg13g2_nor2_2 U1755 (.A(N144), .B(N147), .Y(n395));
sg13g2_nor2_2 U1756 (.A(N199), .B(N202), .Y(n391));
sg13g2_mux2_1 U1757 (.A0(sigma_12), .A1(N316), .S(n1313), .X(n896));
sg13g2_a21oi_2 U1758 (.A1(n398), .A2(kd_12), .B1(N316), .Y(n250));
sg13g2_nor2_2 U1759 (.A(n231), .B(n372), .Y(N324));
sg13g2_inv_2 U1761 (.A(sum_20), .Y(n231));
sg13g2_nor2_2 U1762 (.A(n172), .B(n208), .Y(n252));
sg13g2_mux2_1 U1763 (.A0(sigma_26), .A1(N330), .S(N303), .X(n882));
sg13g2_nor2_2 U1766 (.A(n229), .B(n372), .Y(N325));
sg13g2_nor2_2 U1767 (.A(n229), .B(n381), .Y(N292));
sg13g2_inv_2 U1768 (.A(sum_21), .Y(n229));
sg13g2_inv_2 U1769 (.A(sum_31), .Y(n207));
sg13g2_nor2_2 U1770 (.A(N326), .B(n1307), .Y(n228));
sg13g2_nor2_2 U1771 (.A(n227), .B(n372), .Y(N326));
sg13g2_mux2_1 U1773 (.A0(a_22), .A1(N415), .S(n1296), .X(n851));
sg13g2_nand2_2 U1775 (.A(N559), .B(sum_31), .Y(n562));
sg13g2_nor2_2 U1776 (.A(n225), .B(n372), .Y(N327));
sg13g2_inv_2 U1777 (.A(sum_23), .Y(n225));
sg13g2_inv_2 U1778 (.A(sum_12), .Y(n172));
sg13g2_mux2_1 U1779 (.A0(of_3), .A1(N339), .S(N343), .X(n840));
sg13g2_nor2_2 U1780 (.A(n372), .B(n124), .Y(N313));
sg13g2_inv_2 U1781 (.A(sum_9), .Y(n124));
sg13g2_nor2_2 U1784 (.A(n372), .B(n160), .Y(N319));
sg13g2_inv_2 U1786 (.A(sum_29), .Y(n213));
sg13g2_a21oi_2 U1787 (.A1(product_19), .A2(n292), .B1(n293), .Y(n305));
sg13g2_nor2_2 U1788 (.A(product_23), .B(n293), .Y(n1316));
sg13g2_nor2_2 U1789 (.A(n293), .B(n292), .Y(n1315));
sg13g2_a21oi_2 U1790 (.A1(product_18), .A2(n292), .B1(n293), .Y(n306));
sg13g2_mux2_1 U1791 (.A0(a_30), .A1(N423), .S(net9475), .X(n843));
sg13g2_inv_2 U1792 (.A(n308), .Y(N377));
sg13g2_inv_2 U1793 (.A(n306), .Y(N379));
sg13g2_inv_2 U1795 (.A(n297), .Y(n1308));
sg13g2_mux2_1 U1798 (.A0(p_17), .A1(N378), .S(net9476), .X(n987));
sg13g2_nand3_1 U1799 (.A(n328), .B(n329), .C(n330), .Y(N371));
sg13g2_nand2_2 U1800 (.A(product_10), .B(n292), .Y(n329));
sg13g2_mux2_1 U1801 (.A0(n1312), .A1(n296), .S(net9475), .X(n448));
sg13g2_nor2_2 U1802 (.A(n372), .B(n176), .Y(N315));
sg13g2_inv_2 U1803 (.A(sum_11), .Y(n176));
sg13g2_a21oi_2 U1805 (.A1(product_16), .A2(n292), .B1(n293), .Y(n308));
sg13g2_mux2_1 U1806 (.A0(a_29), .A1(N422), .S(net9476), .X(n844));
sg13g2_mux2_1 U1807 (.A0(n302), .A1(n1328), .S(net14608), .X(n449));
sg13g2_a21oi_2 U1808 (.A1(n292), .A2(product_22), .B1(n293), .Y(n302));
sg13g2_nor2_2 U1810 (.A(state_1_5), .B(state_1_4), .Y(n1298));
sg13g2_mux2_1 U1811 (.A0(n1299), .A1(n305), .S(N360), .X(n450));
sg13g2_o21ai_1 U1813 (.A1(n1301), .A2(n1302), .B1(n1303), .Y(net10403));
sg13g2_inv_2 U1814 (.A(product_26), .Y(n1301));
sg13g2_inv_2 U1815 (.A(n292), .Y(n1302));
sg13g2_inv_2 U1816 (.A(n293), .Y(n1303));
sg13g2_a21oi_2 U1817 (.A1(N263), .A2(sigma_24), .B1(N328), .Y(n224));
sg13g2_inv_2 U1819 (.A(net9475), .Y(net14330));
sg13g2_inv_2 U1820 (.A(net9474), .Y(net9476));
sg13g2_nand4_1 U1821 (.A(n205), .B(n389), .C(n390), .D(n204), .Y(N360));
sg13g2_inv_2 U1822 (.A(n395), .Y(n204));
sg13g2_mux2_1 U1823 (.A0(mr_index_0), .A1(n395), .S(N428), .X(n1007));
sg13g2_mux2_1 U1824 (.A0(md_index_0), .A1(n395), .S(N428), .X(n1005));
sg13g2_nand2_2 U1826 (.A(net11765), .B(n208), .Y(n292));
sg13g2_inv_2 U1828 (.A(state_1_0), .Y(N95));
sg13g2_inv_2 U1829 (.A(net9475), .Y(net14608));
sg13g2_a21oi_2 U1830 (.A1(product_30), .A2(n292), .B1(n293), .Y(n294));
sg13g2_mux2_1 U1831 (.A0(p_24), .A1(net10582), .S(net9475), .X(n980));
sg13g2_a21oi_2 U1833 (.A1(product_24), .A2(n292), .B1(n293), .Y(n300));
sg13g2_inv_2 U1834 (.A(n300), .Y(net10582));
sg13g2_nand3_1 U1835 (.A(n312), .B(n313), .C(n314), .Y(N375));
sg13g2_a21oi_2 U1838 (.A1(sigma_25), .A2(N263), .B1(N329), .Y(n222));
sg13g2_nor2_2 U1839 (.A(n219), .B(n372), .Y(N330));
sg13g2_inv_2 U1840 (.A(sum_26), .Y(n219));
sg13g2_mux2_1 U1841 (.A0(p_12), .A1(N373), .S(net9475), .X(n992));
sg13g2_a21oi_2 U1842 (.A1(product_28), .A2(n292), .B1(n293), .Y(n296));
sg13g2_nor2_2 U1845 (.A(n372), .B(n168), .Y(N317));
sg13g2_inv_2 U1846 (.A(sum_13), .Y(n168));
sg13g2_nand2_2 U1847 (.A(n410), .B(n423), .Y(N136));
sg13g2_nor2_2 U1848 (.A(N263), .B(n396), .Y(n205));
sg13g2_nor2_2 U1849 (.A(n1306), .B(n1314), .Y(n1307));
sg13g2_inv_2 U1851 (.A(sum_8), .Y(n128));
sg13g2_mux2_1 U1852 (.A0(a_12), .A1(N405), .S(net9475), .X(n864));
sg13g2_nor2_2 U1853 (.A(n221), .B(n372), .Y(N329));
sg13g2_a21oi_2 U1855 (.A1(product_27), .A2(n292), .B1(n293), .Y(n297));
sg13g2_inv_2 U1856 (.A(sum_22), .Y(n227));
sg13g2_nor2_2 U1857 (.A(n213), .B(n372), .Y(N333));
sg13g2_mux2_1 U1859 (.A0(a_13), .A1(N406), .S(net9476), .X(n863));
sg13g2_mux2_1 U1861 (.A0(N557), .A1(n291), .S(net9476), .X(n453));
sg13g2_nor2_2 U1862 (.A(n233), .B(n372), .Y(N323));
sg13g2_inv_2 U1863 (.A(sum_19), .Y(n233));
sg13g2_mux2_1 U1864 (.A0(a_8), .A1(N401), .S(net9475), .X(n868));
sg13g2_nor2_2 U1866 (.A(n235), .B(n372), .Y(N322));
sg13g2_mux2_1 U1867 (.A0(p_25), .A1(N386), .S(net9476), .X(n979));
sg13g2_nor2_2 U1869 (.A(n397), .B(N257), .Y(n385));
sg13g2_mux2_1 U1871 (.A0(p_26), .A1(net10403), .S(net9475), .X(n978));
sg13g2_a21oi_2 U1872 (.A1(sigma_30), .A2(N263), .B1(N334), .Y(n212));
sg13g2_inv_2 U1874 (.A(sum_25), .Y(n221));
sg13g2_mux2_1 U1875 (.A0(a_20), .A1(N413), .S(net9475), .X(n853));
sg13g2_mux2_1 U1876 (.A0(a_21), .A1(N414), .S(net9476), .X(n852));
sg13g2_mux2_1 U1877 (.A0(a_18), .A1(N411), .S(net9475), .X(n855));
sg13g2_inv_2 U1878 (.A(sum_18), .Y(n235));
sg13g2_mux2_1 U1880 (.A0(a_24), .A1(N417), .S(net9475), .X(n849));
sg13g2_mux2_1 U1882 (.A0(n1326), .A1(n295), .S(net9476), .X(n454));
sg13g2_nor2_2 U1883 (.A(n164), .B(n208), .Y(n246));
sg13g2_mux2_1 U1885 (.A0(sigma_18), .A1(N322), .S(N303), .X(n890));
sg13g2_nor2_2 U1886 (.A(n217), .B(n372), .Y(N331));
sg13g2_inv_2 U1887 (.A(sum_27), .Y(n217));
sg13g2_mux2_1 U1888 (.A0(N420), .A1(a_27), .S(net13458), .X(n846));
sg13g2_inv_2 U1889 (.A(n303), .Y(n1310));
sg13g2_a21oi_2 U1890 (.A1(product_21), .A2(n292), .B1(n293), .Y(n303));
sg13g2_mux2_1 U1891 (.A0(sigma_22), .A1(N326), .S(n1313), .X(n886));
sg13g2_mux2_1 U1893 (.A0(state_1_1), .A1(N257), .S(N255), .X(n1021));
sg13g2_mux2_1 U1894 (.A0(state_1_7), .A1(N263), .S(N255), .X(n1015));
sg13g2_inv_2 U1895 (.A(N132), .Y(n421));
sg13g2_mux2_1 U1898 (.A0(sigma_28), .A1(N332), .S(N303), .X(n880));
sg13g2_nor2_2 U1899 (.A(n1315), .B(n1316), .Y(N384));
sg13g2_nand2_2 U1900 (.A(n372), .B(n375), .Y(n1313));
sg13g2_nand4_1 U1901 (.A(RS), .B(n399), .C(n35), .D(n36), .Y(n375));
sg13g2_nand2_2 U1903 (.A(n204), .B(n375), .Y(N342));
sg13g2_nand2_2 U1904 (.A(n444), .B(n445), .Y(N180));
sg13g2_nor2_2 U1905 (.A(state_1_4), .B(state_1_3), .Y(n1321));
sg13g2_a21oi_2 U1906 (.A1(product_31), .A2(n292), .B1(n293), .Y(n291));
sg13g2_mux2_1 U1907 (.A0(p_23), .A1(N384), .S(net9476), .X(n981));
sg13g2_nand3_1 U1909 (.A(n1314), .B(n204), .C(n1), .Y(N428));
sg13g2_inv_2 U1910 (.A(n372), .Y(n1317));
sg13g2_nor2_2 U1911 (.A(state_1_2), .B(n1322), .Y(n1323));
sg13g2_nor2_2 U1912 (.A(N161), .B(state_1_1), .Y(n1324));
sg13g2_nor2_2 U1913 (.A(N263), .B(n1317), .Y(net11765));
sg13g2_mux2_1 U1914 (.A0(of_4), .A1(N340), .S(N303), .X(n841));
sg13g2_mux2_1 U1915 (.A0(kpd_13), .A1(sum_13), .S(n397), .X(n959));
sg13g2_mux2_1 U1916 (.A0(kpd_12), .A1(sum_12), .S(n397), .X(n960));
sg13g2_mux2_1 U1917 (.A0(kpd_11), .A1(sum_11), .S(n397), .X(n961));
sg13g2_mux2_1 U1918 (.A0(kpd_10), .A1(sum_10), .S(n397), .X(n962));
sg13g2_mux2_1 U1919 (.A0(kpd_9), .A1(sum_9), .S(n397), .X(n963));
sg13g2_mux2_1 U1920 (.A0(kpd_8), .A1(sum_8), .S(n397), .X(n964));
sg13g2_mux2_1 U1921 (.A0(kpd_7), .A1(sum_7), .S(n397), .X(n965));
sg13g2_mux2_1 U1922 (.A0(kpd_6), .A1(sum_6), .S(n397), .X(n966));
sg13g2_mux2_1 U1923 (.A0(kpd_4), .A1(sum_4), .S(n397), .X(n968));
sg13g2_mux2_1 U1924 (.A0(kpd_5), .A1(sum_5), .S(n397), .X(n967));
sg13g2_mux2_1 U1925 (.A0(kpd_3), .A1(sum_3), .S(n397), .X(n969));
sg13g2_mux2_1 U1926 (.A0(kpd_2), .A1(sum_2), .S(n397), .X(n970));
sg13g2_mux2_1 U1927 (.A0(kpd_1), .A1(sum_1), .S(n397), .X(n971));
sg13g2_mux2_1 U1928 (.A0(kpd_0), .A1(sum_0), .S(n397), .X(n972));
sg13g2_mux2_1 U1929 (.A0(sigma_8), .A1(N312), .S(N303), .X(n900));
sg13g2_mux2_1 U1931 (.A0(a_23), .A1(N416), .S(net9476), .X(n850));
sg13g2_mux2_1 U1932 (.A0(sigma_23), .A1(N327), .S(N303), .X(n885));
sg13g2_nand2_2 U1935 (.A(n373), .B(n374), .Y(N343));
sg13g2_o21ai_1 U1936 (.A1(pv_0), .A2(n206), .B1(n290), .Y(n289));
sg13g2_inv_2 U1939 (.A(n396), .Y(n206));
sg13g2_mux2_1 U1940 (.A0(sigma_25), .A1(N329), .S(N303), .X(n883));
sg13g2_a21oi_2 U1941 (.A1(sigma_16), .A2(N263), .B1(N320), .Y(n240));
sg13g2_nor2_2 U1942 (.A(n223), .B(n372), .Y(N328));
sg13g2_inv_2 U1943 (.A(sum_24), .Y(n223));
sg13g2_inv_2 U1944 (.A(n377), .Y(N340));
sg13g2_inv_2 U1945 (.A(sum_28), .Y(n215));
sg13g2_inv_2 U1946 (.A(sum_30), .Y(n211));
sg13g2_inv_2 U1947 (.A(sum_14), .Y(n164));
sg13g2_mux2_1 U1948 (.A0(a_28), .A1(N421), .S(net9475), .X(n845));
sg13g2_mux2_1 U1949 (.A0(sigma_20), .A1(N324), .S(N303), .X(n888));
sg13g2_mux2_1 U1950 (.A0(sigma_30), .A1(n1241), .S(N303), .X(n878));
sg13g2_inv_2 U1951 (.A(sum_6), .Y(n136));
sg13g2_mux2_1 U1954 (.A0(a_26), .A1(N419), .S(net9475), .X(n847));
sg13g2_nor2_2 U1955 (.A(n237), .B(n372), .Y(N321));
sg13g2_inv_2 U1956 (.A(sum_17), .Y(n237));
sg13g2_mux2_1 U1957 (.A0(kpd_14), .A1(sum_14), .S(n397), .X(n958));
sg13g2_mux2_1 U1959 (.A0(sigma_27), .A1(N331), .S(N303), .X(n881));
sg13g2_mux2_1 U1960 (.A0(a_25), .A1(N418), .S(net9476), .X(n848));
sg13g2_mux2_1 U1961 (.A0(p_16), .A1(N377), .S(net9475), .X(n988));
sg13g2_nor2_2 U1962 (.A(n239), .B(n372), .Y(N320));
sg13g2_inv_2 U1963 (.A(sum_16), .Y(n239));
sg13g2_nor2_2 U1964 (.A(n215), .B(n372), .Y(N332));
sg13g2_nor2_2 U1965 (.A(n211), .B(n372), .Y(N334));
sg13g2_nor2_2 U1967 (.A(N157), .B(N156), .Y(n18));
sg13g2_nor2_2 U1968 (.A(n372), .B(n172), .Y(N316));
sg13g2_nor2_2 U1969 (.A(n372), .B(n180), .Y(N314));
sg13g2_inv_2 U1970 (.A(sum_10), .Y(n180));
sg13g2_mux2_1 U1971 (.A0(a_16), .A1(N409), .S(net9475), .X(n857));
sg13g2_mux2_1 U1972 (.A0(sigma_24), .A1(N328), .S(N303), .X(n884));
sg13g2_mux2_1 U1973 (.A0(kpd_15), .A1(sum_15), .S(n397), .X(n957));
sg13g2_mux2_1 U1974 (.A0(sigma_15), .A1(N319), .S(N303), .X(n893));
sg13g2_nand2_2 U1975 (.A(N552), .B(sum_15), .Y(n558));
sg13g2_mux2_1 U1976 (.A0(a_14), .A1(N407), .S(net9475), .X(n862));
sg13g2_mux2_1 U1977 (.A0(a_15), .A1(N408), .S(net9476), .X(n861));
sg13g2_mux2_1 U1979 (.A0(state_1_9), .A1(n392), .S(N255), .X(n1023));
sg13g2_o21ai_1 U1980 (.A1(n373), .A2(n378), .B1(n377), .Y(N339));
sg13g2_mux2_1 U1982 (.A0(md_index_1), .A1(N430), .S(N428), .X(n1006));
sg13g2_mux2_1 U1983 (.A0(mr_index_1), .A1(N430), .S(N428), .X(n1008));
sg13g2_nor2_2 U1984 (.A(n207), .B(n372), .Y(N335));
sg13g2_inv_2 U1987 (.A(n393), .Y(n372));
sg13g2_mux2_1 U1988 (.A0(state_1_4), .A1(n396), .S(N255), .X(n1018));
sg13g2_nand2_2 U1989 (.A(n372), .B(n375), .Y(N303));
sg13g2_mux2_1 U1990 (.A0(state_1_8), .A1(n393), .S(N255), .X(n1014));
sg13g2_nand2_2 U1991 (.A(n446), .B(N183), .Y(N151));
sg13g2_nand2_2 U1992 (.A(state_1_7), .B(N161), .Y(N174));
sg13g2_mux2_1 U1993 (.A0(state_1_2), .A1(n398), .S(N255), .X(n1020));
sg13g2_mux2_1 U1994 (.A0(state_1_6), .A1(N430), .S(N255), .X(n1016));
sg13g2_nand2_2 U1995 (.A(N128), .B(state_1_2), .Y(N121));
sg13g2_nand2_2 U1996 (.A(state_1_3), .B(N117), .Y(N132));
sg13g2_mux2_1 U1997 (.A0(of_2), .A1(N338), .S(N342), .X(n859));
sg13g2_mux2_1 U1998 (.A0(of_1), .A1(N337), .S(N342), .X(n860));
sg13g2_mux2_1 U1999 (.A0(\err[0][15]), .A1(N359), .S(N342), .X(n941));
sg13g2_mux2_1 U2000 (.A0(\err[0][14]), .A1(N358), .S(N342), .X(n942));
sg13g2_mux2_1 U2001 (.A0(\err[0][13]), .A1(N357), .S(N342), .X(n943));
sg13g2_mux2_1 U2002 (.A0(\err[0][12]), .A1(N356), .S(N342), .X(n944));
sg13g2_mux2_1 U2003 (.A0(\err[0][11]), .A1(N355), .S(N342), .X(n945));
sg13g2_mux2_1 U2004 (.A0(\err[0][10]), .A1(N354), .S(N342), .X(n946));
sg13g2_mux2_1 U2005 (.A0(\err[0][9]), .A1(N353), .S(N342), .X(n947));
sg13g2_mux2_1 U2006 (.A0(\err[0][8]), .A1(N352), .S(N342), .X(n948));
sg13g2_mux2_1 U2007 (.A0(\err[0][7]), .A1(N351), .S(N342), .X(n949));
sg13g2_mux2_1 U2008 (.A0(\err[0][6]), .A1(N350), .S(N342), .X(n950));
sg13g2_mux2_1 U2009 (.A0(\err[0][5]), .A1(N349), .S(N342), .X(n951));
sg13g2_mux2_1 U2010 (.A0(\err[0][0]), .A1(N344), .S(N342), .X(n956));
sg13g2_inv_2 U2012 (.A(n550), .Y(N540));
sg13g2_inv_2 U2013 (.A(N121), .Y(n415));
sg13g2_inv_2 U2015 (.A(n551), .Y(N542));
sg13g2_inv_2 U2016 (.A(i_wb_stb), .Y(N536));
sg13g2_nor2_2 U2057 (.A(\i_wb_data[30]), .B(\i_wb_data[31]), .Y(n1329));
sg13g2_inv_2 U2058 (.A(\i_wb_data[29]), .Y(n463));
sg13g2_inv_2 U2059 (.A(\i_wb_data[28]), .Y(n465));
sg13g2_nor2_2 U2060 (.A(\i_wb_data[27]), .B(N488), .Y(n1330));
sg13g2_inv_2 U2061 (.A(\i_wb_data[25]), .Y(n471));
sg13g2_inv_2 U2062 (.A(\i_wb_data[23]), .Y(n475));
sg13g2_nor2_2 U2063 (.A(\i_wb_data[21]), .B(N494), .Y(n1331));
sg13g2_inv_2 U2064 (.A(\i_wb_data[20]), .Y(n481));
sg13g2_inv_2 U2065 (.A(\i_wb_data[19]), .Y(n483));
sg13g2_nor2_2 U2066 (.A(\i_wb_data[18]), .B(N497), .Y(n1332));
sg13g2_inv_2 U2067 (.A(\i_wb_data[17]), .Y(n487));
sg13g2_inv_2 U2068 (.A(\i_wb_data[16]), .Y(n489));
sg13g2_nor2_2 U2069 (.A(\i_wb_data[15]), .B(N500), .Y(n1333));
sg13g2_inv_2 U2070 (.A(\i_wb_data[14]), .Y(n493));
sg13g2_nor2_2 U2071 (.A(\i_wb_data[12]), .B(N503), .Y(n1334));
sg13g2_inv_2 U2072 (.A(\i_wb_data[11]), .Y(n499));
sg13g2_inv_2 U2073 (.A(\i_wb_data[10]), .Y(n501));
sg13g2_nor2_2 U2074 (.A(\i_wb_adr[14]), .B(\i_wb_adr[15]), .Y(n1335));
sg13g2_nor2_2 U2075 (.A(\i_wb_data[9]), .B(N506), .Y(n1336));
sg13g2_inv_2 U2076 (.A(\i_wb_adr[12]), .Y(n528));
sg13g2_inv_2 U2077 (.A(\i_wb_data[7]), .Y(n507));
sg13g2_nor2_2 U2078 (.A(\i_wb_adr[11]), .B(N525), .Y(n1337));
sg13g2_inv_2 U2079 (.A(\i_wb_adr[10]), .Y(n532));
sg13g2_inv_2 U2080 (.A(\i_wb_data[5]), .Y(n511));
sg13g2_inv_2 U2081 (.A(\i_wb_adr[9]), .Y(n534));
sg13g2_inv_2 U2082 (.A(\i_wb_data[4]), .Y(n513));
sg13g2_nor2_2 U2083 (.A(\i_wb_adr[8]), .B(N528), .Y(n1338));
sg13g2_inv_2 U2084 (.A(\i_wb_adr[7]), .Y(n538));
sg13g2_inv_2 U2085 (.A(i_wb_we), .Y(N534));
sg13g2_xnor2_1 U2086 (.A(N522), .B(\i_wb_adr[3]), .Y(n1345));
sg13g2_xnor2_1 U2087 (.A(\i_wb_adr[2]), .B(\i_wb_adr[5]), .Y(n1344));
sg13g2_inv_2 U2088 (.A(N520), .Y(N521));
sg13g2_inv_2 U2089 (.A(n563), .Y(N559));
sg13g2_inv_2 U2092 (.A(n40), .Y(adr_check));
sg13g2_inv_2 U2093 (.A(\i_wb_data[2]), .Y(n517));
sg13g2_inv_2 U2094 (.A(\i_wb_adr[2]), .Y(n1525));
sg13g2_inv_2 U2095 (.A(\i_wb_adr[6]), .Y(n540));
sg13g2_xnor2_1 U2096 (.A(\i_wb_adr[4]), .B(\i_wb_adr[5]), .Y(n1342));
sg13g2_inv_2 U2097 (.A(n557), .Y(N547));
sg13g2_inv_2 U2098 (.A(n559), .Y(N552));
sg13g2_inv_2 U2101 (.A(\i_wb_adr[3]), .Y(N480));
sg13g2_inv_2 U2102 (.A(\i_wb_adr[4]), .Y(n1341));
sg13g2_inv_2 U2130 (.A(N531), .Y(N532));
sg13g2_inv_2 U2131 (.A(\i_wb_adr[5]), .Y(N522));
sg13g2_nor2_2 U2132 (.A(\i_wb_data[0]), .B(N515), .Y(n1339));
sg13g2_inv_2 U2220 (.A(i_rst), .Y(n1340));
sg13g2_nand2_2 U2221 (.A(N106), .B(state_1_0), .Y(N100));
sg13g2_mux2_1 U2222 (.A0(\o_un[31]), .A1(sigma_31), .S(\i_wb_adr[2]), .X(n1531));
sg13g2_mux2_1 U2223 (.A0(n1348), .A1(n1349), .S(\i_wb_adr[3]), .X(n455));
sg13g2_mux2_1 U2224 (.A0(n1351), .A1(n1352), .S(\i_wb_adr[3]), .X(n458));
sg13g2_mux2_1 U2225 (.A0(n1353), .A1(n1354), .S(\i_wb_adr[5]), .X(n459));
sg13g2_mux2_1 U2226 (.A0(\o_un[30]), .A1(sigma_30), .S(\i_wb_adr[2]), .X(n1532));
sg13g2_mux2_1 U2227 (.A0(n1353), .A1(n1356), .S(\i_wb_adr[5]), .X(n460));
sg13g2_mux2_1 U2228 (.A0(\o_un[29]), .A1(sigma_29), .S(\i_wb_adr[2]), .X(n1533));
sg13g2_mux2_1 U2229 (.A0(n1353), .A1(n1358), .S(\i_wb_adr[5]), .X(n461));
sg13g2_mux2_1 U2230 (.A0(\o_un[28]), .A1(sigma_28), .S(\i_wb_adr[2]), .X(n1534));
sg13g2_mux2_1 U2231 (.A0(n1353), .A1(n1360), .S(\i_wb_adr[5]), .X(n462));
sg13g2_mux2_1 U2232 (.A0(\o_un[27]), .A1(sigma_27), .S(\i_wb_adr[2]), .X(n1535));
sg13g2_mux2_1 U2233 (.A0(n1353), .A1(n1362), .S(\i_wb_adr[5]), .X(n464));
sg13g2_mux2_1 U2234 (.A0(\o_un[26]), .A1(sigma_26), .S(\i_wb_adr[2]), .X(n1536));
sg13g2_mux2_1 U2235 (.A0(n1353), .A1(n1364), .S(\i_wb_adr[5]), .X(n466));
sg13g2_mux2_1 U2236 (.A0(\o_un[25]), .A1(sigma_25), .S(\i_wb_adr[2]), .X(n1537));
sg13g2_mux2_1 U2237 (.A0(n1353), .A1(n1366), .S(\i_wb_adr[5]), .X(n467));
sg13g2_mux2_1 U2238 (.A0(\o_un[24]), .A1(sigma_24), .S(\i_wb_adr[2]), .X(n1538));
sg13g2_mux2_1 U2239 (.A0(n1353), .A1(n1368), .S(\i_wb_adr[5]), .X(n468));
sg13g2_mux2_1 U2240 (.A0(\o_un[23]), .A1(sigma_23), .S(\i_wb_adr[2]), .X(n1539));
sg13g2_mux2_1 U2241 (.A0(n1353), .A1(n1370), .S(\i_wb_adr[5]), .X(n469));
sg13g2_mux2_1 U2242 (.A0(\o_un[22]), .A1(sigma_22), .S(\i_wb_adr[2]), .X(n1540));
sg13g2_mux2_1 U2243 (.A0(n1353), .A1(n1372), .S(\i_wb_adr[5]), .X(n470));
sg13g2_mux2_1 U2244 (.A0(\o_un[21]), .A1(sigma_21), .S(\i_wb_adr[2]), .X(n1541));
sg13g2_mux2_1 U2245 (.A0(n1353), .A1(n1374), .S(\i_wb_adr[5]), .X(n473));
sg13g2_mux2_1 U2246 (.A0(\o_un[20]), .A1(sigma_20), .S(\i_wb_adr[2]), .X(n1542));
sg13g2_mux2_1 U2247 (.A0(n1353), .A1(n1376), .S(\i_wb_adr[5]), .X(n474));
sg13g2_mux2_1 U2248 (.A0(\o_un[19]), .A1(sigma_19), .S(\i_wb_adr[2]), .X(n1543));
sg13g2_mux2_1 U2249 (.A0(n1353), .A1(n1378), .S(\i_wb_adr[5]), .X(n476));
sg13g2_mux2_1 U2250 (.A0(\o_un[18]), .A1(sigma_18), .S(\i_wb_adr[2]), .X(n1544));
sg13g2_mux2_1 U2251 (.A0(n1353), .A1(n1380), .S(\i_wb_adr[5]), .X(n477));
sg13g2_mux2_1 U2252 (.A0(\o_un[17]), .A1(sigma_17), .S(\i_wb_adr[2]), .X(n1545));
sg13g2_mux2_1 U2253 (.A0(n1353), .A1(n1382), .S(\i_wb_adr[5]), .X(n478));
sg13g2_mux2_1 U2254 (.A0(\o_un[16]), .A1(sigma_16), .S(\i_wb_adr[2]), .X(n1546));
sg13g2_mux2_1 U2255 (.A0(n1353), .A1(n1384), .S(\i_wb_adr[5]), .X(n479));
sg13g2_mux2_1 U2256 (.A0(\o_un[15]), .A1(sigma_15), .S(\i_wb_adr[2]), .X(n1547));
sg13g2_mux2_1 U2257 (.A0(n1353), .A1(n1386), .S(\i_wb_adr[5]), .X(n480));
sg13g2_mux2_1 U2258 (.A0(\o_un[14]), .A1(sigma_14), .S(\i_wb_adr[2]), .X(n1548));
sg13g2_mux2_1 U2259 (.A0(n1389), .A1(n1390), .S(\i_wb_adr[3]), .X(n482));
sg13g2_mux2_1 U2260 (.A0(n1392), .A1(n1393), .S(\i_wb_adr[3]), .X(n484));
sg13g2_mux2_1 U2261 (.A0(n1394), .A1(n1395), .S(\i_wb_adr[5]), .X(n485));
sg13g2_mux2_1 U2262 (.A0(\o_un[13]), .A1(sigma_13), .S(\i_wb_adr[2]), .X(n1549));
sg13g2_mux2_1 U2263 (.A0(n1398), .A1(n1399), .S(\i_wb_adr[3]), .X(n486));
sg13g2_mux2_1 U2264 (.A0(n1401), .A1(n1402), .S(\i_wb_adr[3]), .X(n488));
sg13g2_mux2_1 U2265 (.A0(n1403), .A1(n1404), .S(\i_wb_adr[5]), .X(n490));
sg13g2_mux2_1 U2266 (.A0(\o_un[12]), .A1(sigma_12), .S(\i_wb_adr[2]), .X(n1550));
sg13g2_mux2_1 U2267 (.A0(n1407), .A1(n1408), .S(\i_wb_adr[3]), .X(n491));
sg13g2_mux2_1 U2268 (.A0(n1410), .A1(n1411), .S(\i_wb_adr[3]), .X(n492));
sg13g2_mux2_1 U2269 (.A0(n1412), .A1(n1413), .S(\i_wb_adr[5]), .X(n494));
sg13g2_mux2_1 U2270 (.A0(\o_un[11]), .A1(sigma_11), .S(\i_wb_adr[2]), .X(n1551));
sg13g2_mux2_1 U2271 (.A0(n1416), .A1(n1417), .S(\i_wb_adr[3]), .X(n495));
sg13g2_mux2_1 U2272 (.A0(n1419), .A1(n1420), .S(\i_wb_adr[3]), .X(n496));
sg13g2_mux2_1 U2273 (.A0(n1421), .A1(n1422), .S(\i_wb_adr[5]), .X(n497));
sg13g2_mux2_1 U2274 (.A0(\o_un[10]), .A1(sigma_10), .S(\i_wb_adr[2]), .X(n1552));
sg13g2_mux2_1 U2275 (.A0(n1425), .A1(n1426), .S(\i_wb_adr[3]), .X(n498));
sg13g2_mux2_1 U2276 (.A0(n1428), .A1(n1429), .S(\i_wb_adr[3]), .X(n500));
sg13g2_mux2_1 U2277 (.A0(n1430), .A1(n1431), .S(\i_wb_adr[5]), .X(n502));
sg13g2_mux2_1 U2278 (.A0(\o_un[9]), .A1(sigma_9), .S(\i_wb_adr[2]), .X(n1553));
sg13g2_mux2_1 U2279 (.A0(n1434), .A1(n1435), .S(\i_wb_adr[3]), .X(n503));
sg13g2_mux2_1 U2280 (.A0(n1437), .A1(n1438), .S(\i_wb_adr[3]), .X(n504));
sg13g2_mux2_1 U2281 (.A0(n1439), .A1(n1440), .S(\i_wb_adr[5]), .X(n505));
sg13g2_mux2_1 U2282 (.A0(\o_un[8]), .A1(sigma_8), .S(\i_wb_adr[2]), .X(n1554));
sg13g2_mux2_1 U2283 (.A0(n1443), .A1(n1444), .S(\i_wb_adr[3]), .X(n506));
sg13g2_mux2_1 U2284 (.A0(n1446), .A1(n1447), .S(\i_wb_adr[3]), .X(n509));
sg13g2_mux2_1 U2285 (.A0(n1448), .A1(n1449), .S(\i_wb_adr[5]), .X(n510));
sg13g2_mux2_1 U2286 (.A0(\o_un[7]), .A1(sigma_7), .S(\i_wb_adr[2]), .X(n1555));
sg13g2_mux2_1 U2287 (.A0(n1452), .A1(n1453), .S(\i_wb_adr[3]), .X(n512));
sg13g2_mux2_1 U2288 (.A0(n1455), .A1(n1456), .S(\i_wb_adr[3]), .X(n515));
sg13g2_mux2_1 U2289 (.A0(n1457), .A1(n1458), .S(\i_wb_adr[5]), .X(n516));
sg13g2_mux2_1 U2290 (.A0(\o_un[6]), .A1(sigma_6), .S(\i_wb_adr[2]), .X(n1556));
sg13g2_mux2_1 U2291 (.A0(n1461), .A1(n1462), .S(\i_wb_adr[3]), .X(n518));
sg13g2_mux2_1 U2292 (.A0(n1464), .A1(n1465), .S(\i_wb_adr[3]), .X(n519));
sg13g2_mux2_1 U2293 (.A0(n1466), .A1(n1467), .S(\i_wb_adr[5]), .X(n520));
sg13g2_mux2_1 U2294 (.A0(\o_un[5]), .A1(sigma_5), .S(\i_wb_adr[2]), .X(n1557));
sg13g2_mux2_1 U2295 (.A0(n1470), .A1(n1471), .S(\i_wb_adr[3]), .X(n521));
sg13g2_mux2_1 U2296 (.A0(n1473), .A1(n1474), .S(\i_wb_adr[3]), .X(n522));
sg13g2_mux2_1 U2297 (.A0(n1475), .A1(n1476), .S(\i_wb_adr[5]), .X(n523));
sg13g2_mux2_1 U2298 (.A0(\o_un[4]), .A1(sigma_4), .S(\i_wb_adr[2]), .X(n524));
sg13g2_mux2_1 U2299 (.A0(n1479), .A1(n1480), .S(\i_wb_adr[3]), .X(n525));
sg13g2_mux2_1 U2300 (.A0(n1482), .A1(n1483), .S(\i_wb_adr[3]), .X(n526));
sg13g2_mux2_1 U2301 (.A0(n1484), .A1(n1485), .S(\i_wb_adr[5]), .X(n527));
sg13g2_mux2_1 U2302 (.A0(\o_un[3]), .A1(sigma_3), .S(\i_wb_adr[2]), .X(n529));
sg13g2_mux2_1 U2303 (.A0(n1488), .A1(n1489), .S(\i_wb_adr[3]), .X(n530));
sg13g2_mux2_1 U2304 (.A0(n1491), .A1(n1492), .S(\i_wb_adr[3]), .X(n531));
sg13g2_mux2_1 U2305 (.A0(n1493), .A1(n1494), .S(\i_wb_adr[5]), .X(n533));
sg13g2_mux2_1 U2306 (.A0(\o_un[2]), .A1(sigma_2), .S(\i_wb_adr[2]), .X(n535));
sg13g2_mux2_1 U2307 (.A0(n1497), .A1(n1498), .S(\i_wb_adr[3]), .X(n536));
sg13g2_mux2_1 U2308 (.A0(n1500), .A1(n1501), .S(\i_wb_adr[3]), .X(n537));
sg13g2_mux2_1 U2309 (.A0(n1502), .A1(n1503), .S(\i_wb_adr[5]), .X(n539));
sg13g2_mux2_1 U2310 (.A0(\o_un[1]), .A1(sigma_1), .S(\i_wb_adr[2]), .X(n541));
sg13g2_mux2_1 U2311 (.A0(n1506), .A1(n1507), .S(\i_wb_adr[3]), .X(n543));
sg13g2_mux2_1 U2312 (.A0(n1509), .A1(n1510), .S(\i_wb_adr[3]), .X(n544));
sg13g2_mux2_1 U2313 (.A0(n1511), .A1(n1512), .S(\i_wb_adr[5]), .X(n545));
sg13g2_mux2_1 U2314 (.A0(\o_un[0]), .A1(sigma_0), .S(\i_wb_adr[2]), .X(n546));
sg13g2_mux2_1 U2315 (.A0(n1515), .A1(n1516), .S(\i_wb_adr[3]), .X(n547));
sg13g2_mux2_1 U2316 (.A0(n1518), .A1(n1519), .S(\i_wb_adr[3]), .X(n548));
sg13g2_mux2_1 U2317 (.A0(n1520), .A1(n1521), .S(\i_wb_adr[5]), .X(n552));
sg13g2_nor2_2 U2318 (.A(n1344), .B(n1522), .Y(n1523));
sg13g2_mux2_1 U2319 (.A0(n1523), .A1(rl_6), .S(n1345), .X(n553));
sg13g2_nand2_2 U2320 (.A(of_0), .B(n1525), .Y(n1524));
sg13g2_nand2_2 U2321 (.A(of_1), .B(n1525), .Y(n1526));
sg13g2_nand2_2 U2322 (.A(of_2), .B(n1525), .Y(n1527));
sg13g2_nand2_2 U2323 (.A(of_3), .B(n1525), .Y(n1528));
sg13g2_nand2_2 U2324 (.A(of_4), .B(n1525), .Y(n1529));
sg13g2_mux2_1 U2325 (.A0(\err[0][15]), .A1(\err[1][15]), .S(\i_wb_adr[2]), .X(n554));
sg13g2_mux2_1 U2326 (.A0(pv_15), .A1(kpd_15), .S(\i_wb_adr[2]), .X(n555));
sg13g2_mux2_1 U2327 (.A0(kd_15), .A1(sp_15), .S(\i_wb_adr[2]), .X(n556));
sg13g2_mux2_1 U2328 (.A0(kp_15), .A1(ki_15), .S(\i_wb_adr[2]), .X(n561));
sg13g2_mux2_1 U2329 (.A0(n1350), .A1(n1347), .S(\i_wb_adr[4]), .X(n564));
sg13g2_nand2_2 U2330 (.A(n1531), .B(n1530), .Y(n1354));
sg13g2_nand2_2 U2331 (.A(n1532), .B(n1530), .Y(n1356));
sg13g2_nand2_2 U2332 (.A(n1533), .B(n1530), .Y(n1358));
sg13g2_nand2_2 U2333 (.A(n1534), .B(n1530), .Y(n1360));
sg13g2_nand2_2 U2334 (.A(n1535), .B(n1530), .Y(n1362));
sg13g2_nand2_2 U2335 (.A(n1536), .B(n1530), .Y(n1364));
sg13g2_nand2_2 U2336 (.A(n1537), .B(n1530), .Y(n1366));
sg13g2_nand2_2 U2337 (.A(n1538), .B(n1530), .Y(n1368));
sg13g2_nand2_2 U2338 (.A(n1539), .B(n1530), .Y(n1370));
sg13g2_nand2_2 U2339 (.A(n1540), .B(n1530), .Y(n1372));
sg13g2_nand2_2 U2340 (.A(n1541), .B(n1530), .Y(n1374));
sg13g2_nand2_2 U2341 (.A(n1542), .B(n1530), .Y(n1376));
sg13g2_nand2_2 U2342 (.A(n1543), .B(n1530), .Y(n1378));
sg13g2_nand2_2 U2343 (.A(n1544), .B(n1530), .Y(n1380));
sg13g2_nand2_2 U2344 (.A(n1545), .B(n1530), .Y(n1382));
sg13g2_nand2_2 U2345 (.A(n1546), .B(n1530), .Y(n1384));
sg13g2_nand2_2 U2346 (.A(n1547), .B(n1530), .Y(n1386));
sg13g2_mux2_1 U2347 (.A0(\err[0][14]), .A1(\err[1][14]), .S(\i_wb_adr[2]), .X(n565));
sg13g2_mux2_1 U2348 (.A0(pv_14), .A1(kpd_14), .S(\i_wb_adr[2]), .X(n566));
sg13g2_mux2_1 U2349 (.A0(kd_14), .A1(sp_14), .S(\i_wb_adr[2]), .X(n567));
sg13g2_mux2_1 U2350 (.A0(kp_14), .A1(ki_14), .S(\i_wb_adr[2]), .X(n571));
sg13g2_mux2_1 U2351 (.A0(n1391), .A1(n1388), .S(\i_wb_adr[4]), .X(n572));
sg13g2_nand2_2 U2352 (.A(n1548), .B(n1530), .Y(n1395));
sg13g2_mux2_1 U2353 (.A0(\err[0][13]), .A1(\err[1][13]), .S(\i_wb_adr[2]), .X(n573));
sg13g2_mux2_1 U2354 (.A0(pv_13), .A1(kpd_13), .S(\i_wb_adr[2]), .X(n574));
sg13g2_mux2_1 U2355 (.A0(kd_13), .A1(sp_13), .S(\i_wb_adr[2]), .X(n575));
sg13g2_mux2_1 U2356 (.A0(kp_13), .A1(ki_13), .S(\i_wb_adr[2]), .X(n576));
sg13g2_mux2_1 U2357 (.A0(n1400), .A1(n1397), .S(\i_wb_adr[4]), .X(n577));
sg13g2_nand2_2 U2358 (.A(n1549), .B(n1530), .Y(n1404));
sg13g2_mux2_1 U2359 (.A0(\err[0][12]), .A1(\err[1][12]), .S(\i_wb_adr[2]), .X(n578));
sg13g2_mux2_1 U2360 (.A0(pv_12), .A1(kpd_12), .S(\i_wb_adr[2]), .X(n579));
sg13g2_mux2_1 U2361 (.A0(kd_12), .A1(sp_12), .S(\i_wb_adr[2]), .X(n580));
sg13g2_mux2_1 U2362 (.A0(kp_12), .A1(ki_12), .S(\i_wb_adr[2]), .X(n581));
sg13g2_mux2_1 U2363 (.A0(n1409), .A1(n1406), .S(\i_wb_adr[4]), .X(n582));
sg13g2_nand2_2 U2364 (.A(n1550), .B(n1530), .Y(n1413));
sg13g2_mux2_1 U2365 (.A0(\err[0][11]), .A1(\err[1][11]), .S(\i_wb_adr[2]), .X(n583));
sg13g2_mux2_1 U2366 (.A0(pv_11), .A1(kpd_11), .S(\i_wb_adr[2]), .X(n584));
sg13g2_mux2_1 U2367 (.A0(kd_11), .A1(sp_11), .S(\i_wb_adr[2]), .X(n585));
sg13g2_mux2_1 U2368 (.A0(kp_11), .A1(ki_11), .S(\i_wb_adr[2]), .X(n586));
sg13g2_mux2_1 U2369 (.A0(n1418), .A1(n1415), .S(\i_wb_adr[4]), .X(n587));
sg13g2_nand2_2 U2370 (.A(n1551), .B(n1530), .Y(n1422));
sg13g2_mux2_1 U2371 (.A0(\err[0][10]), .A1(\err[1][10]), .S(\i_wb_adr[2]), .X(n588));
sg13g2_mux2_1 U2372 (.A0(pv_10), .A1(kpd_10), .S(\i_wb_adr[2]), .X(n589));
sg13g2_mux2_1 U2373 (.A0(kd_10), .A1(sp_10), .S(\i_wb_adr[2]), .X(n590));
sg13g2_mux2_1 U2374 (.A0(kp_10), .A1(ki_10), .S(\i_wb_adr[2]), .X(n591));
sg13g2_mux2_1 U2375 (.A0(n1427), .A1(n1424), .S(\i_wb_adr[4]), .X(n592));
sg13g2_nand2_2 U2376 (.A(n1552), .B(n1530), .Y(n1431));
sg13g2_mux2_1 U2377 (.A0(\err[0][9]), .A1(\err[1][9]), .S(\i_wb_adr[2]), .X(n593));
sg13g2_mux2_1 U2378 (.A0(pv_9), .A1(kpd_9), .S(\i_wb_adr[2]), .X(n594));
sg13g2_mux2_1 U2379 (.A0(kd_9), .A1(sp_9), .S(\i_wb_adr[2]), .X(n595));
sg13g2_mux2_1 U2380 (.A0(kp_9), .A1(ki_9), .S(\i_wb_adr[2]), .X(n596));
sg13g2_mux2_1 U2381 (.A0(n1436), .A1(n1433), .S(\i_wb_adr[4]), .X(n597));
sg13g2_nand2_2 U2382 (.A(n1553), .B(n1530), .Y(n1440));
sg13g2_mux2_1 U2383 (.A0(\err[0][8]), .A1(\err[1][8]), .S(\i_wb_adr[2]), .X(n598));
sg13g2_mux2_1 U2384 (.A0(pv_8), .A1(kpd_8), .S(\i_wb_adr[2]), .X(n599));
sg13g2_mux2_1 U2385 (.A0(kd_8), .A1(sp_8), .S(\i_wb_adr[2]), .X(n600));
sg13g2_mux2_1 U2386 (.A0(kp_8), .A1(ki_8), .S(\i_wb_adr[2]), .X(n601));
sg13g2_mux2_1 U2387 (.A0(n1445), .A1(n1442), .S(\i_wb_adr[4]), .X(n602));
sg13g2_nand2_2 U2388 (.A(n1554), .B(n1530), .Y(n1449));
sg13g2_mux2_1 U2389 (.A0(\err[0][7]), .A1(\err[1][7]), .S(\i_wb_adr[2]), .X(n603));
sg13g2_mux2_1 U2390 (.A0(pv_7), .A1(kpd_7), .S(\i_wb_adr[2]), .X(n604));
sg13g2_mux2_1 U2391 (.A0(kd_7), .A1(sp_7), .S(\i_wb_adr[2]), .X(n605));
sg13g2_mux2_1 U2392 (.A0(kp_7), .A1(ki_7), .S(\i_wb_adr[2]), .X(n606));
sg13g2_mux2_1 U2393 (.A0(n1454), .A1(n1451), .S(\i_wb_adr[4]), .X(n607));
sg13g2_nand2_2 U2394 (.A(n1555), .B(n1530), .Y(n1458));
sg13g2_mux2_1 U2395 (.A0(\err[0][6]), .A1(\err[1][6]), .S(\i_wb_adr[2]), .X(n608));
sg13g2_mux2_1 U2396 (.A0(pv_6), .A1(kpd_6), .S(\i_wb_adr[2]), .X(n609));
sg13g2_mux2_1 U2397 (.A0(kd_6), .A1(sp_6), .S(\i_wb_adr[2]), .X(n610));
sg13g2_mux2_1 U2398 (.A0(kp_6), .A1(ki_6), .S(\i_wb_adr[2]), .X(n611));
sg13g2_mux2_1 U2399 (.A0(n1463), .A1(n1460), .S(\i_wb_adr[4]), .X(n612));
sg13g2_nand2_2 U2400 (.A(n1556), .B(n1530), .Y(n1467));
sg13g2_mux2_1 U2401 (.A0(\err[0][5]), .A1(\err[1][5]), .S(\i_wb_adr[2]), .X(n613));
sg13g2_mux2_1 U2402 (.A0(pv_5), .A1(kpd_5), .S(\i_wb_adr[2]), .X(n614));
sg13g2_mux2_1 U2403 (.A0(kd_5), .A1(sp_5), .S(\i_wb_adr[2]), .X(n615));
sg13g2_mux2_1 U2404 (.A0(kp_5), .A1(ki_5), .S(\i_wb_adr[2]), .X(n616));
sg13g2_mux2_1 U2405 (.A0(n1472), .A1(n1469), .S(\i_wb_adr[4]), .X(n617));
sg13g2_nand2_2 U2406 (.A(n1557), .B(n1530), .Y(n1476));
sg13g2_mux2_1 U2407 (.A0(n1477), .A1(n1529), .S(\i_wb_adr[3]), .X(n618));
sg13g2_mux2_1 U2408 (.A0(\err[0][4]), .A1(\err[1][4]), .S(\i_wb_adr[2]), .X(n619));
sg13g2_mux2_1 U2409 (.A0(pv_4), .A1(kpd_4), .S(\i_wb_adr[2]), .X(n620));
sg13g2_mux2_1 U2410 (.A0(kd_4), .A1(sp_4), .S(\i_wb_adr[2]), .X(n621));
sg13g2_mux2_1 U2411 (.A0(kp_4), .A1(ki_4), .S(\i_wb_adr[2]), .X(n622));
sg13g2_mux2_1 U2412 (.A0(n1481), .A1(n1478), .S(\i_wb_adr[4]), .X(n623));
sg13g2_nand2_2 U2413 (.A(n1558), .B(n1341), .Y(n1485));
sg13g2_mux2_1 U2414 (.A0(n1486), .A1(n1528), .S(\i_wb_adr[3]), .X(n624));
sg13g2_mux2_1 U2415 (.A0(\err[0][3]), .A1(\err[1][3]), .S(\i_wb_adr[2]), .X(n625));
sg13g2_mux2_1 U2416 (.A0(pv_3), .A1(kpd_3), .S(\i_wb_adr[2]), .X(n626));
sg13g2_mux2_1 U2417 (.A0(kd_3), .A1(sp_3), .S(\i_wb_adr[2]), .X(n627));
sg13g2_mux2_1 U2418 (.A0(kp_3), .A1(ki_3), .S(\i_wb_adr[2]), .X(n628));
sg13g2_mux2_1 U2419 (.A0(n1490), .A1(n1487), .S(\i_wb_adr[4]), .X(n629));
sg13g2_nand2_2 U2420 (.A(n1559), .B(n1341), .Y(n1494));
sg13g2_mux2_1 U2421 (.A0(n1495), .A1(n1527), .S(\i_wb_adr[3]), .X(n630));
sg13g2_mux2_1 U2422 (.A0(\err[0][2]), .A1(\err[1][2]), .S(\i_wb_adr[2]), .X(n631));
sg13g2_mux2_1 U2423 (.A0(pv_2), .A1(kpd_2), .S(\i_wb_adr[2]), .X(n632));
sg13g2_mux2_1 U2424 (.A0(kd_2), .A1(sp_2), .S(\i_wb_adr[2]), .X(n633));
sg13g2_mux2_1 U2425 (.A0(kp_2), .A1(ki_2), .S(\i_wb_adr[2]), .X(n634));
sg13g2_mux2_1 U2426 (.A0(n1499), .A1(n1496), .S(\i_wb_adr[4]), .X(n635));
sg13g2_nand2_2 U2427 (.A(n1560), .B(n1341), .Y(n1503));
sg13g2_mux2_1 U2428 (.A0(n1504), .A1(n1526), .S(\i_wb_adr[3]), .X(n636));
sg13g2_mux2_1 U2429 (.A0(\err[0][1]), .A1(\err[1][1]), .S(\i_wb_adr[2]), .X(n637));
sg13g2_mux2_1 U2430 (.A0(pv_1), .A1(kpd_1), .S(\i_wb_adr[2]), .X(n638));
sg13g2_mux2_1 U2431 (.A0(kd_1), .A1(sp_1), .S(\i_wb_adr[2]), .X(n639));
sg13g2_mux2_1 U2432 (.A0(kp_1), .A1(ki_1), .S(\i_wb_adr[2]), .X(n640));
sg13g2_mux2_1 U2433 (.A0(n1508), .A1(n1505), .S(\i_wb_adr[4]), .X(n641));
sg13g2_nand2_2 U2434 (.A(n1561), .B(n1341), .Y(n1512));
sg13g2_mux2_1 U2435 (.A0(n1513), .A1(n1524), .S(\i_wb_adr[3]), .X(n642));
sg13g2_mux2_1 U2436 (.A0(\err[0][0]), .A1(\err[1][0]), .S(\i_wb_adr[2]), .X(n643));
sg13g2_mux2_1 U2437 (.A0(pv_0), .A1(kpd_0), .S(\i_wb_adr[2]), .X(n644));
sg13g2_mux2_1 U2438 (.A0(kd_0), .A1(sp_0), .S(\i_wb_adr[2]), .X(n645));
sg13g2_mux2_1 U2439 (.A0(kp_0), .A1(ki_0), .S(\i_wb_adr[2]), .X(n646));
sg13g2_mux2_1 U2440 (.A0(n1517), .A1(n1514), .S(\i_wb_adr[4]), .X(n647));
sg13g2_nand2_2 U2441 (.A(n1562), .B(n1341), .Y(n1521));
sg13g2_nor2_2 U2442 (.A(n1563), .B(n1564), .Y(N39));
sg13g2_mux2_1 U2443 (.A0(n1565), .A1(n1341), .S(\i_wb_adr[3]), .X(n648));
sg13g2_mux2_1 U2444 (.A0(n1341), .A1(n1525), .S(\i_wb_adr[3]), .X(n649));
sg13g2_mux2_1 U2445 (.A0(\wl[0]), .A1(wl_3), .S(n1566), .X(n650));
sg13g2_o21ai_1 U2446 (.A1(\i_wb_adr[4]), .A2(n542), .B1(\i_wb_adr[2]), .Y(n1565));
sg13g2_dfrbp_2 wack_reg (.CLK(i_clk), .D(n1105), .Q(wack), .Q_N(N537), .RESET_B(n1340));
sg13g2_dfrbp_1 wla_reg (.CLK(i_clk), .D(n1106), .Q(\wl[0]), .Q_N(n542), .RESET_B(n1340));
sg13g2_dfrbp_1 wlb_reg (.CLK(i_clk), .D(n1010), .Q(wl_3), .RESET_B(n1340));
adder_32bit_0 adder_32bit_0(.\i_a[0](a_0), .\i_a[1](a_1), .\i_a[2](a_2), .\i_a[3](a_3), .\i_a[4](a_4), .\i_a[5](a_5), .\i_a[6](a_6), .\i_a[7](a_7), .\i_a[8](a_8), .\i_a[9](a_9), .\i_a[10](a_10), .\i_a[11](a_11), .\i_a[12](a_12), .\i_a[13](a_13), .\i_a[14](a_14), .\i_a[15](a_15), .\i_a[16](a_16), .\i_a[17](a_17), .\i_a[18](a_18), .\i_a[19](a_19), .\i_a[20](a_20), .\i_a[21](a_21), .\i_a[22](a_22), .\i_a[23](a_23), .\i_a[24](a_24), .\i_a[25](a_25), .\i_a[26](a_26), .\i_a[27](a_27), .\i_a[28](a_28), .\i_a[29](a_29), .\i_a[30](a_30), .\i_a[31](a_31), .\i_b[0](p_0), .\i_b[1](p_1), .\i_b[2](p_2), .\i_b[3](p_3), .\i_b[4](p_4), .\i_b[5](p_5), .\i_b[6](p_6), .\i_b[7](p_7), .\i_b[8](p_8), .\i_b[9](p_9), .\i_b[10](p_10), .\i_b[11](p_11), .\i_b[12](p_12), .\i_b[13](p_13), .\i_b[14](p_14), .\i_b[15](p_15), .\i_b[16](p_16), .\i_b[17](p_17), .\i_b[18](p_18), .\i_b[19](p_19), .\i_b[20](p_20), .\i_b[21](p_21), .\i_b[22](p_22), .\i_b[23](p_23), .\i_b[24](p_24), .\i_b[25](p_25), .\i_b[26](p_26), .\i_b[27](p_27), .\i_b[28](p_28), .\i_b[29](p_29), .\i_b[30](p_30), .\i_b[31](p_31), .\o_s[0](sum_0), .\o_s[1](sum_1), .\o_s[2](sum_2), .\o_s[3](sum_3), .\o_s[4](sum_4), .\o_s[5](sum_5), .\o_s[6](sum_6), .\o_s[7](sum_7), .\o_s[8](sum_8), .\o_s[9](sum_9), .\o_s[10](sum_10), .\o_s[11](sum_11), .\o_s[12](sum_12), .\o_s[13](sum_13), .\o_s[14](sum_14), .\o_s[15](sum_15), .\o_s[16](sum_16), .\o_s[17](sum_17), .\o_s[18](sum_18), .\o_s[19](sum_19), .\o_s[20](sum_20), .\o_s[21](sum_21), .\o_s[22](sum_22), .\o_s[23](sum_23), .\o_s[24](sum_24), .\o_s[25](sum_25), .\o_s[26](sum_26), .\o_s[27](sum_27), .\o_s[28](sum_28), .\o_s[29](sum_29), .\o_s[30](sum_30), .\o_s[31](sum_31), .i_c(cout), .o_c());
multiplier_16x16bit_pipelined multiplier_16x16bit_pipelined(.\i_md[0](md_0), .\i_md[1](md_1), .\i_md[2](md_2), .\i_md[3](md_3), .\i_md[4](md_4), .\i_md[5](md_5), .\i_md[6](md_6), .\i_md[7](md_7), .\i_md[8](md_8), .\i_md[9](md_9), .\i_md[10](md_10), .\i_md[11](md_11), .\i_md[12](md_12), .\i_md[13](md_13), .\i_md[14](md_14), .\i_md[15](md_15), .\i_mr[0](mr_0), .\i_mr[1](mr_1), .\i_mr[2](mr_2), .\i_mr[3](mr_3), .\i_mr[4](mr_4), .\i_mr[5](mr_5), .\i_mr[6](mr_6), .\i_mr[7](mr_7), .\i_mr[8](mr_8), .\i_mr[9](mr_9), .\i_mr[10](mr_10), .\i_mr[11](mr_11), .\i_mr[12](mr_12), .\i_mr[13](mr_13), .\i_mr[14](mr_14), .\i_mr[15](mr_15), .\o_product[0](product_0), .\o_product[1](product_1), .\o_product[2](product_2), .\o_product[3](product_3), .\o_product[4](product_4), .\o_product[5](product_5), .\o_product[6](product_6), .\o_product[7](product_7), .\o_product[8](product_8), .\o_product[9](product_9), .\o_product[10](product_10), .\o_product[11](product_11), .\o_product[12](product_12), .\o_product[13](product_13), .\o_product[14](product_14), .\o_product[15](product_15), .\o_product[16](product_16), .\o_product[17](product_17), .\o_product[18](product_18), .\o_product[19](product_19), .\o_product[20](product_20), .\o_product[21](product_21), .\o_product[22](product_22), .\o_product[23](product_23), .\o_product[24](product_24), .\o_product[25](product_25), .\o_product[26](product_26), .\o_product[27](product_27), .\o_product[28](product_28), .\o_product[29](product_29), .\o_product[30](product_30), .\o_product[31](product_31), .i_clk(i_clk), .i_rst(n1340), .i_start(start), .o_ready());
endmodule

module adder_32bit_0 (\i_a[0], \i_a[1], \i_a[2], \i_a[3], \i_a[4], \i_a[5], \i_a[6], \i_a[7], \i_a[8], \i_a[9], \i_a[10], \i_a[11], \i_a[12], \i_a[13], \i_a[14], \i_a[15], \i_a[16], \i_a[17], \i_a[18], \i_a[19], \i_a[20], \i_a[21], \i_a[22], \i_a[23], \i_a[24], \i_a[25], \i_a[26], \i_a[27], \i_a[28], \i_a[29], \i_a[30], \i_a[31], \i_b[0], \i_b[1], \i_b[2], \i_b[3], \i_b[4], \i_b[5], \i_b[6], \i_b[7], \i_b[8], \i_b[9], \i_b[10], \i_b[11], \i_b[12], \i_b[13], \i_b[14], \i_b[15], \i_b[16], \i_b[17], \i_b[18], \i_b[19], \i_b[20], \i_b[21], \i_b[22], \i_b[23], \i_b[24], \i_b[25], \i_b[26], \i_b[27], \i_b[28], \i_b[29], \i_b[30], \i_b[31], \o_s[0], \o_s[1], \o_s[2], \o_s[3], \o_s[4], \o_s[5], \o_s[6], \o_s[7], \o_s[8], \o_s[9], \o_s[10], \o_s[11], \o_s[12], \o_s[13], \o_s[14], \o_s[15], \o_s[16], \o_s[17], \o_s[18], \o_s[19], \o_s[20], \o_s[21], \o_s[22], \o_s[23], \o_s[24], \o_s[25], \o_s[26], \o_s[27], \o_s[28], \o_s[29], \o_s[30], \o_s[31], i_c, o_c);
input \i_a[0], \i_a[1], \i_a[2], \i_a[3], \i_a[4], \i_a[5], \i_a[6], \i_a[7], \i_a[8], \i_a[9], \i_a[10], \i_a[11], \i_a[12], \i_a[13], \i_a[14], \i_a[15], \i_a[16], \i_a[17], \i_a[18], \i_a[19], \i_a[20], \i_a[21], \i_a[22], \i_a[23], \i_a[24], \i_a[25], \i_a[26], \i_a[27], \i_a[28], \i_a[29], \i_a[30], \i_a[31], \i_b[0], \i_b[1], \i_b[2], \i_b[3], \i_b[4], \i_b[5], \i_b[6], \i_b[7], \i_b[8], \i_b[9], \i_b[10], \i_b[11], \i_b[12], \i_b[13], \i_b[14], \i_b[15], \i_b[16], \i_b[17], \i_b[18], \i_b[19], \i_b[20], \i_b[21], \i_b[22], \i_b[23], \i_b[24], \i_b[25], \i_b[26], \i_b[27], \i_b[28], \i_b[29], \i_b[30], \i_b[31], i_c;
output \o_s[0], \o_s[1], \o_s[2], \o_s[3], \o_s[4], \o_s[5], \o_s[6], \o_s[7], \o_s[8], \o_s[9], \o_s[10], \o_s[11], \o_s[12], \o_s[13], \o_s[14], \o_s[15], \o_s[16], \o_s[17], \o_s[18], \o_s[19], \o_s[20], \o_s[21], \o_s[22], \o_s[23], \o_s[24], \o_s[25], \o_s[26], \o_s[27], \o_s[28], \o_s[29], \o_s[30], \o_s[31], o_c;

sg13g2_inv_2 U1 (.A(n1), .Y(\o_s[9]));
sg13g2_xnor2_1 U2 (.A(P0_9), .B(G4_4), .Y(n1));
sg13g2_inv_2 U3 (.A(n14), .Y(\o_s[26]));
sg13g2_xnor2_1 U4 (.A(P0_8), .B(G6_7), .Y(n2));
sg13g2_inv_2 U5 (.A(n3), .Y(\o_s[7]));
sg13g2_xnor2_1 U6 (.A(P0_7), .B(G3_3), .Y(n3));
sg13g2_inv_2 U7 (.A(n13), .Y(\o_s[27]));
sg13g2_xnor2_1 U8 (.A(P0_6), .B(G6_5), .Y(n4));
sg13g2_inv_2 U9 (.A(n5), .Y(\o_s[5]));
sg13g2_xnor2_1 U10 (.A(P0_5), .B(G3_2), .Y(n5));
sg13g2_inv_2 U11 (.A(n6), .Y(\o_s[4]));
sg13g2_xnor2_1 U12 (.A(P0_4), .B(G6_3), .Y(n6));
sg13g2_inv_2 U13 (.A(n7), .Y(\o_s[3]));
sg13g2_xnor2_1 U14 (.A(P0_3), .B(G2_1), .Y(n7));
sg13g2_xnor2_1 U15 (.A(P0_27), .B(G5_13), .Y(n13));
sg13g2_inv_2 U16 (.A(n27), .Y(\o_s[14]));
sg13g2_xnor2_1 U17 (.A(P0_14), .B(G6_13), .Y(n27));
sg13g2_xnor2_1 U18 (.A(P0_15), .B(G4_7), .Y(n26));
sg13g2_inv_2 U19 (.A(n10), .Y(\o_s[2]));
sg13g2_xnor2_1 U20 (.A(P0_2), .B(G6_1), .Y(n10));
sg13g2_inv_2 U21 (.A(P0_31), .Y(n35));
sg13g2_xnor2_1 U22 (.A(P0_20), .B(G6_19), .Y(n20));
sg13g2_o21ai_1 U23 (.A1(G6_15), .A2(P0_16), .B1(n36), .Y(n25));
sg13g2_xnor2_1 U24 (.A(n35), .B(G5_15), .Y(\o_s[31]));
sg13g2_inv_2 U25 (.A(n12), .Y(\o_s[28]));
sg13g2_xnor2_1 U26 (.A(P0_30), .B(\G6[29]), .Y(n9));
sg13g2_xnor2_1 U27 (.A(P0_12), .B(G6_11), .Y(n29));
sg13g2_inv_2 U28 (.A(n19), .Y(\o_s[21]));
sg13g2_inv_2 U29 (.A(n15), .Y(\o_s[25]));
sg13g2_xnor2_1 U30 (.A(P0_25), .B(G5_12), .Y(n15));
sg13g2_xnor2_1 U31 (.A(P0_21), .B(G5_10), .Y(n19));
sg13g2_xnor2_1 U32 (.A(P0_24), .B(G6_23), .Y(n16));
sg13g2_inv_2 U33 (.A(n17), .Y(\o_s[23]));
sg13g2_xnor2_1 U34 (.A(P0_23), .B(G5_11), .Y(n17));
sg13g2_inv_2 U35 (.A(G1_0), .Y(n8));
sg13g2_inv_2 U36 (.A(n8), .Y(n33));
sg13g2_inv_2 U37 (.A(n11), .Y(\o_s[29]));
sg13g2_xnor2_1 U38 (.A(G5_14), .B(P0_29), .Y(n11));
sg13g2_inv_2 U39 (.A(n20), .Y(\o_s[20]));
sg13g2_nand2_2 U40 (.A(G6_15), .B(P0_16), .Y(n36));
sg13g2_inv_2 U41 (.A(n21), .Y(\o_s[1]));
sg13g2_xnor2_1 U42 (.A(n38), .B(n33), .Y(n21));
sg13g2_inv_2 U43 (.A(n22), .Y(\o_s[19]));
sg13g2_xnor2_1 U44 (.A(P0_19), .B(G5_9), .Y(n22));
sg13g2_inv_2 U45 (.A(n25), .Y(\o_s[16]));
sg13g2_inv_2 U46 (.A(n23), .Y(\o_s[18]));
sg13g2_inv_2 U47 (.A(n24), .Y(\o_s[17]));
sg13g2_xnor2_1 U48 (.A(P0_17), .B(G5_8), .Y(n24));
sg13g2_inv_2 U49 (.A(n2), .Y(\o_s[8]));
sg13g2_inv_2 U50 (.A(n29), .Y(\o_s[12]));
sg13g2_inv_2 U51 (.A(n26), .Y(\o_s[15]));
sg13g2_xnor2_1 U52 (.A(P0_22), .B(G6_21), .Y(n18));
sg13g2_xnor2_1 U53 (.A(P0_28), .B(G6_27), .Y(n12));
sg13g2_inv_2 U54 (.A(n16), .Y(\o_s[24]));
sg13g2_inv_2 U55 (.A(n28), .Y(\o_s[13]));
sg13g2_xnor2_1 U56 (.A(P0_13), .B(G4_6), .Y(n28));
sg13g2_xnor2_1 U57 (.A(P0_26), .B(G6_25), .Y(n14));
sg13g2_inv_2 U58 (.A(n9), .Y(\o_s[30]));
sg13g2_inv_2 U59 (.A(n30), .Y(\o_s[11]));
sg13g2_xnor2_1 U60 (.A(P0_11), .B(G4_5), .Y(n30));
sg13g2_xnor2_1 U61 (.A(P0_18), .B(G6_17), .Y(n23));
sg13g2_inv_2 U62 (.A(n31), .Y(\o_s[10]));
sg13g2_inv_2 U63 (.A(n32), .Y(\o_s[0]));
sg13g2_xnor2_1 U64 (.A(i_c), .B(P0_0), .Y(n32));
sg13g2_xnor2_1 U65 (.A(P0_10), .B(G6_9), .Y(n31));
sg13g2_inv_2 U66 (.A(P0_1), .Y(n37));
sg13g2_inv_2 U67 (.A(n37), .Y(n38));
sg13g2_inv_2 U68 (.A(n4), .Y(\o_s[6]));
sg13g2_inv_2 U69 (.A(n18), .Y(\o_s[22]));
operator_A_0 operator_A_0(.A(\i_a[0]), .B(\i_b[0]), .G(G0_0), .P(P0_0));
operator_A_33 operator_A_31(.A(\i_a[31]), .B(\i_b[31]), .G(G0_31), .P(P0_31));
operator_A_34 operator_A_30(.A(\i_a[30]), .B(\i_b[30]), .G(G0_30), .P(P0_30));
operator_A_35 operator_A_29(.A(\i_a[29]), .B(\i_b[29]), .G(G0_29), .P(P0_29));
operator_A_36 operator_A_28(.A(\i_a[28]), .B(\i_b[28]), .G(G0_28), .P(P0_28));
operator_A_37 operator_A_27(.A(\i_a[27]), .B(\i_b[27]), .G(G0_27), .P(P0_27));
operator_A_38 operator_A_26(.A(\i_a[26]), .B(\i_b[26]), .G(G0_26), .P(P0_26));
operator_A_39 operator_A_25(.A(\i_a[25]), .B(\i_b[25]), .G(G0_25), .P(P0_25));
operator_A_40 operator_A_24(.A(\i_a[24]), .B(\i_b[24]), .G(G0_24), .P(P0_24));
operator_A_41 operator_A_23(.A(\i_a[23]), .B(\i_b[23]), .G(G0_23), .P(P0_23));
operator_A_42 operator_A_22(.A(\i_a[22]), .B(\i_b[22]), .G(G0_22), .P(P0_22));
operator_A_43 operator_A_21(.A(\i_a[21]), .B(\i_b[21]), .G(G0_21), .P(P0_21));
operator_A_44 operator_A_20(.A(\i_a[20]), .B(\i_b[20]), .G(G0_20), .P(P0_20));
operator_A_45 operator_A_19(.A(\i_a[19]), .B(\i_b[19]), .G(G0_19), .P(P0_19));
operator_A_46 operator_A_18(.A(\i_a[18]), .B(\i_b[18]), .G(G0_18), .P(P0_18));
operator_A_47 operator_A_17(.A(\i_a[17]), .B(\i_b[17]), .G(G0_17), .P(P0_17));
operator_A_48 operator_A_16(.A(\i_a[16]), .B(\i_b[16]), .G(G0_16), .P(P0_16));
operator_A_49 operator_A_15(.A(\i_a[15]), .B(\i_b[15]), .G(G0_15), .P(P0_15));
operator_A_50 operator_A_14(.A(\i_a[14]), .B(\i_b[14]), .G(G0_14), .P(P0_14));
operator_A_51 operator_A_13(.A(\i_a[13]), .B(\i_b[13]), .G(G0_13), .P(P0_13));
operator_A_52 operator_A_12(.A(\i_a[12]), .B(\i_b[12]), .G(G0_12), .P(P0_12));
operator_A_53 operator_A_11(.A(\i_a[11]), .B(\i_b[11]), .G(G0_11), .P(P0_11));
operator_A_54 operator_A_10(.A(\i_a[10]), .B(\i_b[10]), .G(G0_10), .P(P0_10));
operator_A_55 operator_A_9(.A(\i_a[9]), .B(\i_b[9]), .G(G0_9), .P(P0_9));
operator_A_56 operator_A_8(.A(\i_a[8]), .B(\i_b[8]), .G(G0_8), .P(P0_8));
operator_A_57 operator_A_7(.A(\i_a[7]), .B(\i_b[7]), .G(G0_7), .P(P0_7));
operator_A_58 operator_A_6(.A(\i_a[6]), .B(\i_b[6]), .G(G0_6), .P(P0_6));
operator_A_59 operator_A_5(.A(\i_a[5]), .B(\i_b[5]), .G(G0_5), .P(P0_5));
operator_A_60 operator_A_4(.A(\i_a[4]), .B(\i_b[4]), .G(G0_4), .P(P0_4));
operator_A_61 operator_A_3(.A(\i_a[3]), .B(\i_b[3]), .G(G0_3), .P(P0_3));
operator_A_62 operator_A_2(.A(\i_a[2]), .B(\i_b[2]), .G(G0_2), .P(P0_2));
operator_A_63 operator_A_1(.A(\i_a[1]), .B(\i_b[1]), .G(G0_1), .P(P0_1));
operator_B_0 operator_B_stage_1_1(.G(G0_2), .G1(G0_1), .Go(G1_1), .P(P0_2), .P1(P0_1), .Po(P1_1));
operator_B_50 operator_B_stage_4_15(.G(G3_15), .G1(G3_11), .Go(G4_15), .P(P3_15), .P1(P3_11), .Po(P4_15));
operator_B_51 operator_B_stage_4_14(.G(G3_14), .G1(G3_10), .Go(G4_14), .P(P3_14), .P1(P3_10), .Po(P4_14));
operator_B_52 operator_B_stage_4_13(.G(G3_13), .G1(G3_9), .Go(G4_13), .P(P3_13), .P1(P3_9), .Po(P4_13));
operator_B_53 operator_B_stage_4_12(.G(G3_12), .G1(G3_8), .Go(G4_12), .P(P3_12), .P1(P3_8), .Po(P4_12));
operator_B_54 operator_B_stage_4_11(.G(G3_11), .G1(G3_7), .Go(G4_11), .P(P3_11), .P1(P3_7), .Po(P4_11));
operator_B_55 operator_B_stage_4_10(.G(G3_10), .G1(G3_6), .Go(G4_10), .P(P3_10), .P1(P3_6), .Po(P4_10));
operator_B_56 operator_B_stage_4_9(.G(G3_9), .G1(G3_5), .Go(G4_9), .P(P3_9), .P1(P3_5), .Po(P4_9));
operator_B_57 operator_B_stage_4_8(.G(G3_8), .G1(G3_4), .Go(G4_8), .P(P3_8), .P1(P3_4), .Po(P4_8));
operator_B_58 operator_B_stage_3_15(.G(G2_15), .G1(G2_13), .Go(G3_15), .P(P2_15), .P1(P2_13), .Po(P3_15));
operator_B_59 operator_B_stage_3_14(.G(G2_14), .G1(G2_12), .Go(G3_14), .P(P2_14), .P1(P2_12), .Po(P3_14));
operator_B_60 operator_B_stage_3_13(.G(G2_13), .G1(G2_11), .Go(G3_13), .P(P2_13), .P1(P2_11), .Po(P3_13));
operator_B_61 operator_B_stage_3_12(.G(G2_12), .G1(G2_10), .Go(G3_12), .P(P2_12), .P1(P2_10), .Po(P3_12));
operator_B_62 operator_B_stage_3_11(.G(G2_11), .G1(G2_9), .Go(G3_11), .P(P2_11), .P1(P2_9), .Po(P3_11));
operator_B_63 operator_B_stage_3_10(.G(G2_10), .G1(G2_8), .Go(G3_10), .P(P2_10), .P1(P2_8), .Po(P3_10));
operator_B_64 operator_B_stage_3_9(.G(G2_9), .G1(G2_7), .Go(G3_9), .P(P2_9), .P1(P2_7), .Po(P3_9));
operator_B_65 operator_B_stage_3_8(.G(G2_8), .G1(G2_6), .Go(G3_8), .P(P2_8), .P1(P2_6), .Po(P3_8));
operator_B_66 operator_B_stage_3_7(.G(G2_7), .G1(G2_5), .Go(G3_7), .P(P2_7), .P1(P2_5), .Po(P3_7));
operator_B_67 operator_B_stage_3_6(.G(G2_6), .G1(G2_4), .Go(G3_6), .P(P2_6), .P1(P2_4), .Po(P3_6));
operator_B_68 operator_B_stage_3_5(.G(G2_5), .G1(G2_3), .Go(G3_5), .P(P2_5), .P1(P2_3), .Po(P3_5));
operator_B_69 operator_B_stage_3_4(.G(G2_4), .G1(G2_2), .Go(G3_4), .P(P2_4), .P1(P2_2), .Po(P3_4));
operator_B_70 operator_B_stage_2_15(.G(G1_15), .G1(G1_14), .Go(G2_15), .P(P1_15), .P1(P1_14), .Po(P2_15));
operator_B_71 operator_B_stage_2_14(.G(G1_14), .G1(G1_13), .Go(G2_14), .P(P1_14), .P1(P1_13), .Po(P2_14));
operator_B_72 operator_B_stage_2_13(.G(G1_13), .G1(G1_12), .Go(G2_13), .P(P1_13), .P1(P1_12), .Po(P2_13));
operator_B_73 operator_B_stage_2_12(.G(G1_12), .G1(G1_11), .Go(G2_12), .P(P1_12), .P1(P1_11), .Po(P2_12));
operator_B_74 operator_B_stage_2_11(.G(G1_11), .G1(G1_10), .Go(G2_11), .P(P1_11), .P1(P1_10), .Po(P2_11));
operator_B_75 operator_B_stage_2_10(.G(G1_10), .G1(G1_9), .Go(G2_10), .P(P1_10), .P1(P1_9), .Po(P2_10));
operator_B_76 operator_B_stage_2_9(.G(G1_9), .G1(G1_8), .Go(G2_9), .P(P1_9), .P1(P1_8), .Po(P2_9));
operator_B_77 operator_B_stage_2_8(.G(G1_8), .G1(G1_7), .Go(G2_8), .P(P1_8), .P1(P1_7), .Po(P2_8));
operator_B_78 operator_B_stage_2_7(.G(G1_7), .G1(G1_6), .Go(G2_7), .P(P1_7), .P1(P1_6), .Po(P2_7));
operator_B_79 operator_B_stage_2_6(.G(G1_6), .G1(G1_5), .Go(G2_6), .P(P1_6), .P1(P1_5), .Po(P2_6));
operator_B_80 operator_B_stage_2_5(.G(G1_5), .G1(G1_4), .Go(G2_5), .P(P1_5), .P1(P1_4), .Po(P2_5));
operator_B_81 operator_B_stage_2_4(.G(G1_4), .G1(G1_3), .Go(G2_4), .P(P1_4), .P1(P1_3), .Po(P2_4));
operator_B_82 operator_B_stage_2_3(.G(G1_3), .G1(G1_2), .Go(G2_3), .P(P1_3), .P1(P1_2), .Po(P2_3));
operator_B_83 operator_B_stage_2_2(.G(G1_2), .G1(G1_1), .Go(G2_2), .P(P1_2), .P1(P1_1), .Po(P2_2));
operator_B_84 operator_B_stage_1_15(.G(G0_30), .G1(G0_29), .Go(G1_15), .P(P0_30), .P1(P0_29), .Po(P1_15));
operator_B_85 operator_B_stage_1_14(.G(G0_28), .G1(G0_27), .Go(G1_14), .P(P0_28), .P1(P0_27), .Po(P1_14));
operator_B_86 operator_B_stage_1_13(.G(G0_26), .G1(G0_25), .Go(G1_13), .P(P0_26), .P1(P0_25), .Po(P1_13));
operator_B_87 operator_B_stage_1_12(.G(G0_24), .G1(G0_23), .Go(G1_12), .P(P0_24), .P1(P0_23), .Po(P1_12));
operator_B_88 operator_B_stage_1_11(.G(G0_22), .G1(G0_21), .Go(G1_11), .P(P0_22), .P1(P0_21), .Po(P1_11));
operator_B_89 operator_B_stage_1_10(.G(G0_20), .G1(G0_19), .Go(G1_10), .P(P0_20), .P1(P0_19), .Po(P1_10));
operator_B_90 operator_B_stage_1_9(.G(G0_18), .G1(G0_17), .Go(G1_9), .P(P0_18), .P1(P0_17), .Po(P1_9));
operator_B_91 operator_B_stage_1_8(.G(G0_16), .G1(G0_15), .Go(G1_8), .P(P0_16), .P1(P0_15), .Po(P1_8));
operator_B_92 operator_B_stage_1_7(.G(G0_14), .G1(G0_13), .Go(G1_7), .P(P0_14), .P1(P0_13), .Po(P1_7));
operator_B_93 operator_B_stage_1_6(.G(G0_12), .G1(G0_11), .Go(G1_6), .P(P0_12), .P1(P0_11), .Po(P1_6));
operator_B_94 operator_B_stage_1_5(.G(G0_10), .G1(G0_9), .Go(G1_5), .P(P0_10), .P1(P0_9), .Po(P1_5));
operator_B_95 operator_B_stage_1_4(.G(G0_8), .G1(G0_7), .Go(G1_4), .P(P0_8), .P1(P0_7), .Po(P1_4));
operator_B_96 operator_B_stage_1_3(.G(G0_6), .G1(G0_5), .Go(G1_3), .P(P0_6), .P1(P0_5), .Po(P1_3));
operator_B_97 operator_B_stage_1_2(.G(G0_4), .G1(G0_3), .Go(G1_2), .P(P0_4), .P1(P0_3), .Po(P1_2));
operator_C_0 operator_C_stage_1_0(.G(G0_0), .G1(i_c), .Go(G1_0), .P(P0_0));
operator_C_33 operator_C_stage_6_15(.G(G0_31), .G1(G5_15), .Go(o_c), .P(P0_31));
operator_C_34 operator_C_stage_6_14(.G(G0_29), .G1(G5_14), .Go(\G6[29]), .P(P0_29));
operator_C_35 operator_C_stage_6_13(.G(G0_27), .G1(G5_13), .Go(G6_27), .P(P0_27));
operator_C_36 operator_C_stage_6_12(.G(G0_25), .G1(G5_12), .Go(G6_25), .P(P0_25));
operator_C_37 operator_C_stage_6_11(.G(G0_23), .G1(G5_11), .Go(G6_23), .P(P0_23));
operator_C_38 operator_C_stage_6_10(.G(G0_21), .G1(G5_10), .Go(G6_21), .P(P0_21));
operator_C_39 operator_C_stage_6_9(.G(G0_19), .G1(G5_9), .Go(G6_19), .P(P0_19));
operator_C_40 operator_C_stage_6_8(.G(G0_17), .G1(G5_8), .Go(G6_17), .P(P0_17));
operator_C_41 operator_C_stage_6_7(.G(G0_15), .G1(G4_7), .Go(G6_15), .P(P0_15));
operator_C_42 operator_C_stage_6_6(.G(G0_13), .G1(G4_6), .Go(G6_13), .P(P0_13));
operator_C_43 operator_C_stage_6_5(.G(G0_11), .G1(G4_5), .Go(G6_11), .P(P0_11));
operator_C_44 operator_C_stage_6_4(.G(G0_9), .G1(G4_4), .Go(G6_9), .P(P0_9));
operator_C_45 operator_C_stage_6_3(.G(G0_7), .G1(G3_3), .Go(G6_7), .P(P0_7));
operator_C_46 operator_C_stage_6_2(.G(G0_5), .G1(G3_2), .Go(G6_5), .P(P0_5));
operator_C_47 operator_C_stage_6_1(.G(G0_3), .G1(G2_1), .Go(G6_3), .P(P0_3));
operator_C_48 operator_C_stage_6_0(.G(G0_1), .G1(G1_0), .Go(G6_1), .P(n38));
operator_C_49 operator_C_stage_5_15(.G(G4_15), .G1(G4_7), .Go(G5_15), .P(P4_15));
operator_C_50 operator_C_stage_5_14(.G(G4_14), .G1(G4_6), .Go(G5_14), .P(P4_14));
operator_C_51 operator_C_stage_5_13(.G(G4_13), .G1(G4_5), .Go(G5_13), .P(P4_13));
operator_C_52 operator_C_stage_5_12(.G(G4_12), .G1(G4_4), .Go(G5_12), .P(P4_12));
operator_C_53 operator_C_stage_5_11(.G(G4_11), .G1(G3_3), .Go(G5_11), .P(P4_11));
operator_C_54 operator_C_stage_5_10(.G(G4_10), .G1(G3_2), .Go(G5_10), .P(P4_10));
operator_C_55 operator_C_stage_5_9(.G(G4_9), .G1(G2_1), .Go(G5_9), .P(P4_9));
operator_C_56 operator_C_stage_5_8(.G(G4_8), .G1(n33), .Go(G5_8), .P(P4_8));
operator_C_57 operator_C_stage_4_7(.G(G3_7), .G1(G3_3), .Go(G4_7), .P(P3_7));
operator_C_58 operator_C_stage_4_6(.G(G3_6), .G1(G3_2), .Go(G4_6), .P(P3_6));
operator_C_59 operator_C_stage_4_5(.G(G3_5), .G1(G2_1), .Go(G4_5), .P(P3_5));
operator_C_60 operator_C_stage_4_4(.G(G3_4), .G1(n33), .Go(G4_4), .P(P3_4));
operator_C_61 operator_C_stage_3_3(.G(G2_3), .G1(G2_1), .Go(G3_3), .P(P2_3));
operator_C_62 operator_C_stage_3_2(.G(G2_2), .G1(G1_0), .Go(G3_2), .P(P2_2));
operator_C_63 operator_C_stage_2_1(.G(G1_1), .G1(G1_0), .Go(G2_1), .P(P1_1));
endmodule

module operator_A_0 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n1), .Y(P));
sg13g2_inv_2 U2 (.A(n2), .Y(G));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n1));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n2));
endmodule

module operator_A_33 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_34 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(A), .B(B), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(P));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_35 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_36 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_37 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_38 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_39 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_40 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_41 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_42 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_43 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(P));
sg13g2_xnor2_1 U4 (.A(A), .B(B), .Y(n4));
endmodule

module operator_A_44 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_45 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_46 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(A), .Y(n3));
sg13g2_nand2_2 U2 (.A(n5), .B(n6), .Y(n8));
sg13g2_inv_2 U3 (.A(n7), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n7));
sg13g2_nand2_2 U5 (.A(A), .B(B), .Y(n5));
sg13g2_nand2_2 U6 (.A(n3), .B(n4), .Y(n6));
sg13g2_inv_2 U7 (.A(B), .Y(n4));
sg13g2_inv_2 U8 (.A(n8), .Y(P));
endmodule

module operator_A_47 (A, B, G, P);
input A, B;
output G, P;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(G));
sg13g2_inv_2 U3 (.A(n4), .Y(P));
sg13g2_xnor2_1 U4 (.A(A), .B(B), .Y(n4));
endmodule

module operator_A_48 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_49 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_50 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_51 (A, B, G, P);
input A, B;
output G, P;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(G));
sg13g2_inv_2 U3 (.A(n4), .Y(P));
sg13g2_xnor2_1 U4 (.A(A), .B(B), .Y(n4));
endmodule

module operator_A_52 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_53 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_54 (A, B, G, P);
input A, B;
output G, P;

sg13g2_o21ai_1 U1 (.A1(A), .A2(B), .B1(n3), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(P));
sg13g2_inv_2 U3 (.A(n4), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n4));
sg13g2_nand2_2 U5 (.A(A), .B(B), .Y(n3));
endmodule

module operator_A_55 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(P));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_56 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_57 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_58 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_59 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_60 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_inv_2 U2 (.A(n3), .Y(G));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_61 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_62 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_63 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_B_0 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(Po));
sg13g2_inv_2 U3 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_B_50 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_51 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_52 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_53 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_54 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_55 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_56 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_57 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_58 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_59 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_60 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_61 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_62 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n5), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n5));
sg13g2_inv_2 U3 (.A(n4), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n4));
endmodule

module operator_B_63 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Go));
sg13g2_nor2_2 U2 (.A(n1), .B(n3), .Y(Po));
sg13g2_inv_2 U3 (.A(P1), .Y(n1));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n4));
sg13g2_inv_2 U5 (.A(P), .Y(n3));
endmodule

module operator_B_64 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_65 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_66 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_67 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_68 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_69 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_70 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_71 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_72 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_73 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_74 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_75 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n4));
sg13g2_inv_2 U3 (.A(n5), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n5));
endmodule

module operator_B_76 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_77 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_78 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U3 (.A(n1), .Y(Po));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_79 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(Po));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_80 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_81 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_82 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_83 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_84 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_85 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_86 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_87 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_88 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_89 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_90 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P), .B(P1), .Y(n4));
endmodule

module operator_B_91 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_92 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_93 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n4));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n5));
sg13g2_inv_2 U4 (.A(n5), .Y(Po));
endmodule

module operator_B_94 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_95 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_96 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_97 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_C_0 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(Go));
endmodule

module operator_C_33 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_34 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_35 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_36 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_37 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_38 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_39 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_40 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_41 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n3));
endmodule

module operator_C_42 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n3));
endmodule

module operator_C_43 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_44 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_45 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_46 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_47 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_48 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_49 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_50 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_51 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_52 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_53 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_54 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n5), .Y(Go));
sg13g2_nor2_2 U2 (.A(n4), .B(G), .Y(n5));
sg13g2_nor2_2 U3 (.A(n2), .B(n3), .Y(n4));
sg13g2_inv_2 U4 (.A(P), .Y(n2));
sg13g2_inv_2 U5 (.A(G1), .Y(n3));
endmodule

module operator_C_55 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_56 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_57 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_58 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_59 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(G1), .Y(n3));
sg13g2_nor2_2 U2 (.A(n4), .B(G), .Y(n5));
sg13g2_inv_2 U3 (.A(n5), .Y(Go));
sg13g2_nor2_2 U4 (.A(n2), .B(n3), .Y(n4));
sg13g2_inv_2 U5 (.A(P), .Y(n2));
endmodule

module operator_C_60 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_61 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_62 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_63 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module multiplier_16x16bit_pipelined (\i_md[0], \i_md[1], \i_md[2], \i_md[3], \i_md[4], \i_md[5], \i_md[6], \i_md[7], \i_md[8], \i_md[9], \i_md[10], \i_md[11], \i_md[12], \i_md[13], \i_md[14], \i_md[15], \i_mr[0], \i_mr[1], \i_mr[2], \i_mr[3], \i_mr[4], \i_mr[5], \i_mr[6], \i_mr[7], \i_mr[8], \i_mr[9], \i_mr[10], \i_mr[11], \i_mr[12], \i_mr[13], \i_mr[14], \i_mr[15], \o_product[0], \o_product[1], \o_product[2], \o_product[3], \o_product[4], \o_product[5], \o_product[6], \o_product[7], \o_product[8], \o_product[9], \o_product[10], \o_product[11], \o_product[12], \o_product[13], \o_product[14], \o_product[15], \o_product[16], \o_product[17], \o_product[18], \o_product[19], \o_product[20], \o_product[21], \o_product[22], \o_product[23], \o_product[24], \o_product[25], \o_product[26], \o_product[27], \o_product[28], \o_product[29], \o_product[30], \o_product[31], i_clk, i_rst, i_start, o_ready);
input \i_md[0], \i_md[1], \i_md[2], \i_md[3], \i_md[4], \i_md[5], \i_md[6], \i_md[7], \i_md[8], \i_md[9], \i_md[10], \i_md[11], \i_md[12], \i_md[13], \i_md[14], \i_md[15], \i_mr[0], \i_mr[1], \i_mr[2], \i_mr[3], \i_mr[4], \i_mr[5], \i_mr[6], \i_mr[7], \i_mr[8], \i_mr[9], \i_mr[10], \i_mr[11], \i_mr[12], \i_mr[13], \i_mr[14], \i_mr[15], i_clk, i_rst, i_start;
output \o_product[0], \o_product[1], \o_product[2], \o_product[3], \o_product[4], \o_product[5], \o_product[6], \o_product[7], \o_product[8], \o_product[9], \o_product[10], \o_product[11], \o_product[12], \o_product[13], \o_product[14], \o_product[15], \o_product[16], \o_product[17], \o_product[18], \o_product[19], \o_product[20], \o_product[21], \o_product[22], \o_product[23], \o_product[24], \o_product[25], \o_product[26], \o_product[27], \o_product[28], \o_product[29], \o_product[30], \o_product[31], o_ready;

sg13g2_dfrbp_2 \md_reg[0] (.CLK(i_clk), .D(n314), .Q(md_0), .Q_N(n93), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[1] (.CLK(i_clk), .D(n315), .Q(md_1), .Q_N(n95), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[2] (.CLK(i_clk), .D(n316), .Q(md_2), .Q_N(n97), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[3] (.CLK(i_clk), .D(n317), .Q(md_3), .Q_N(n99), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[4] (.CLK(i_clk), .D(n318), .Q(md_4), .Q_N(n101), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[5] (.CLK(i_clk), .D(n319), .Q(md_5), .Q_N(n103), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[6] (.CLK(i_clk), .D(n320), .Q(md_6), .Q_N(n105), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[7] (.CLK(i_clk), .D(n321), .Q(md_7), .Q_N(n107), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[8] (.CLK(i_clk), .D(n322), .Q(md_8), .Q_N(n109), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[9] (.CLK(i_clk), .D(n323), .Q(md_9), .Q_N(n111), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[10] (.CLK(i_clk), .D(n324), .Q(md_10), .Q_N(n113), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[11] (.CLK(i_clk), .D(n325), .Q(md_11), .Q_N(n115), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[12] (.CLK(i_clk), .D(n326), .Q(md_12), .Q_N(n117), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[13] (.CLK(i_clk), .D(n327), .Q(md_13), .Q_N(n119), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[14] (.CLK(i_clk), .D(n328), .Q(md_14), .Q_N(n121), .RESET_B(i_rst));
sg13g2_dfrbp_2 \md_reg[15] (.CLK(i_clk), .D(n329), .Q(md_15), .Q_N(n123), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[0] (.CLK(i_clk), .D(n298), .Q(mr_0), .Q_N(n61), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[1] (.CLK(i_clk), .D(n299), .Q(mr_1), .Q_N(n63), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[2] (.CLK(i_clk), .D(n300), .Q(mr_2), .Q_N(n65), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[3] (.CLK(i_clk), .D(n301), .Q(mr_3), .Q_N(n67), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[4] (.CLK(i_clk), .D(n302), .Q(mr_4), .Q_N(n69), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[5] (.CLK(i_clk), .D(n303), .Q(mr_5), .Q_N(n71), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[6] (.CLK(i_clk), .D(n304), .Q(mr_6), .Q_N(n73), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[7] (.CLK(i_clk), .D(n305), .Q(mr_7), .Q_N(n75), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[8] (.CLK(i_clk), .D(n306), .Q(mr_8), .Q_N(n77), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[9] (.CLK(i_clk), .D(n307), .Q(mr_9), .Q_N(n79), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[10] (.CLK(i_clk), .D(n308), .Q(mr_10), .Q_N(n81), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[11] (.CLK(i_clk), .D(n309), .Q(mr_11), .Q_N(n83), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[12] (.CLK(i_clk), .D(n310), .Q(mr_12), .Q_N(n85), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[13] (.CLK(i_clk), .D(n311), .Q(mr_13), .Q_N(n87), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[14] (.CLK(i_clk), .D(n312), .Q(mr_14), .Q_N(n89), .RESET_B(i_rst));
sg13g2_dfrbp_2 \mr_reg[15] (.CLK(i_clk), .D(n313), .Q(mr_15), .Q_N(n91), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w0_reg[0] (.CLK(i_clk), .D(n291), .Q(reg_layer_2_w0_0), .Q_N(n49), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w0_reg[1] (.CLK(i_clk), .D(n292), .Q(reg_layer_2_w0_1), .Q_N(n51), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w2_reg[0] (.CLK(i_clk), .D(n287), .Q(reg_layer_2_w2_0), .Q_N(n41), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w2_reg[1] (.CLK(i_clk), .D(n288), .Q(reg_layer_2_w2_1), .Q_N(n43), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w2_reg[2] (.CLK(i_clk), .D(n289), .Q(reg_layer_2_w2_2), .Q_N(n45), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w3_reg[0] (.CLK(i_clk), .D(n285), .Q(reg_layer_2_w3_0), .Q_N(n37), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w3_reg[1] (.CLK(i_clk), .D(n286), .Q(reg_layer_2_w3_1), .Q_N(n39), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w4_reg[0] (.CLK(i_clk), .D(n283), .Q(reg_layer_2_w4_0), .Q_N(n33), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w4_reg[1] (.CLK(i_clk), .D(n284), .Q(reg_layer_2_w4_1), .Q_N(n35), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w5_reg[0] (.CLK(i_clk), .D(n281), .Q(reg_layer_2_w5_0), .Q_N(n29), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w5_reg[1] (.CLK(i_clk), .D(n282), .Q(reg_layer_2_w5_1), .Q_N(n31), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w6_reg[0] (.CLK(i_clk), .D(n279), .Q(reg_layer_2_w6_0), .Q_N(n25), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w6_reg[1] (.CLK(i_clk), .D(n280), .Q(reg_layer_2_w6_1), .Q_N(n27), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w7_reg[0] (.CLK(i_clk), .D(n277), .Q(reg_layer_2_w7_0), .Q_N(n21), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w7_reg[1] (.CLK(i_clk), .D(n278), .Q(reg_layer_2_w7_1), .Q_N(n23), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w8_reg[0] (.CLK(i_clk), .D(n275), .Q(reg_layer_2_w8_0), .Q_N(n17), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w8_reg[1] (.CLK(i_clk), .D(n276), .Q(reg_layer_2_w8_1), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w9_reg[0] (.CLK(i_clk), .D(n273), .Q(reg_layer_2_w9_0), .Q_N(n13), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w9_reg[1] (.CLK(i_clk), .D(n274), .Q(reg_layer_2_w9_1), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w10_reg[0] (.CLK(i_clk), .D(n271), .Q(reg_layer_2_w10_0), .Q_N(n9), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w10_reg[1] (.CLK(i_clk), .D(n272), .Q(reg_layer_2_w10_1), .Q_N(n11), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w11_reg[0] (.CLK(i_clk), .D(n267), .Q(reg_layer_2_w11_0), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w11_reg[1] (.CLK(i_clk), .D(n268), .Q(reg_layer_2_w11_1), .Q_N(n3), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w11_reg[2] (.CLK(i_clk), .D(n269), .Q(reg_layer_2_w11_2), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w11_reg[3] (.CLK(i_clk), .D(n270), .Q(reg_layer_2_w11_3), .Q_N(n7), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w12_reg[0] (.CLK(i_clk), .D(n264), .Q(reg_layer_2_w12_0), .Q_N(n213), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w12_reg[1] (.CLK(i_clk), .D(n265), .Q(reg_layer_2_w12_1), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w12_reg[2] (.CLK(i_clk), .D(n266), .Q(reg_layer_2_w12_2), .Q_N(n217), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w13_reg[0] (.CLK(i_clk), .D(n261), .Q(reg_layer_2_w13_0), .Q_N(n207), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w13_reg[1] (.CLK(i_clk), .D(n262), .Q(reg_layer_2_w13_1), .Q_N(n209), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w13_reg[2] (.CLK(i_clk), .D(n263), .Q(reg_layer_2_w13_2), .Q_N(n211), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w14_reg[0] (.CLK(i_clk), .D(n258), .Q(reg_layer_2_w14_0), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w14_reg[1] (.CLK(i_clk), .D(n259), .Q(reg_layer_2_w14_1), .Q_N(n203), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w14_reg[2] (.CLK(i_clk), .D(n260), .Q(reg_layer_2_w14_2), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w15_reg[0] (.CLK(i_clk), .D(n255), .Q(reg_layer_2_w15_0), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w15_reg[1] (.CLK(i_clk), .D(n256), .Q(reg_layer_2_w15_1), .Q_N(n197), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w15_reg[2] (.CLK(i_clk), .D(n257), .Q(reg_layer_2_w15_2), .Q_N(n199), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w16_reg[0] (.CLK(i_clk), .D(n251), .Q(reg_layer_2_w16_0), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w16_reg[1] (.CLK(i_clk), .D(n252), .Q(reg_layer_2_w16_1), .Q_N(n190), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w16_reg[2] (.CLK(i_clk), .D(n253), .Q(reg_layer_2_w16_2), .Q_N(n192), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w16_reg[3] (.CLK(i_clk), .D(n254), .Q(reg_layer_2_w16_3), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w17_reg[0] (.CLK(i_clk), .D(n248), .Q(reg_layer_2_w17_0), .Q_N(n182), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w17_reg[1] (.CLK(i_clk), .D(n249), .Q(reg_layer_2_w17_1), .Q_N(n184), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w17_reg[2] (.CLK(i_clk), .D(n250), .Q(reg_layer_2_w17_2), .Q_N(n186), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w18_reg[0] (.CLK(i_clk), .D(n244), .Q(reg_layer_2_w18_0), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w18_reg[1] (.CLK(i_clk), .D(n245), .Q(reg_layer_2_w18_1), .Q_N(n176), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w18_reg[2] (.CLK(i_clk), .D(n246), .Q(reg_layer_2_w18_2), .Q_N(n178), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w18_reg[3] (.CLK(i_clk), .D(n247), .Q(reg_layer_2_w18_3), .Q_N(n180), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w19_reg[0] (.CLK(i_clk), .D(n241), .Q(reg_layer_2_w19_0), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w19_reg[1] (.CLK(i_clk), .D(n242), .Q(reg_layer_2_w19_1), .Q_N(n170), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w19_reg[2] (.CLK(i_clk), .D(n243), .Q(reg_layer_2_w19_2), .Q_N(n172), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w20_reg[0] (.CLK(i_clk), .D(n237), .Q(reg_layer_2_w20_0), .Q_N(n160), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w20_reg[1] (.CLK(i_clk), .D(n238), .Q(reg_layer_2_w20_1), .Q_N(n162), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w20_reg[2] (.CLK(i_clk), .D(n239), .Q(reg_layer_2_w20_2), .Q_N(n164), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w20_reg[3] (.CLK(i_clk), .D(n240), .Q(reg_layer_2_w20_3), .Q_N(n166), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w21_reg[0] (.CLK(i_clk), .D(n234), .Q(reg_layer_2_w21_0), .Q_N(n155), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w21_reg[1] (.CLK(i_clk), .D(n235), .Q(reg_layer_2_w21_1), .Q_N(n157), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w21_reg[2] (.CLK(i_clk), .D(n236), .Q(reg_layer_2_w21_2), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w22_reg[0] (.CLK(i_clk), .D(n232), .Q(reg_layer_2_w22_0), .Q_N(n151), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w22_reg[1] (.CLK(i_clk), .D(n233), .Q(reg_layer_2_w22_1), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w23_reg[0] (.CLK(i_clk), .D(n230), .Q(reg_layer_2_w23_0), .Q_N(n147), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w23_reg[1] (.CLK(i_clk), .D(n231), .Q(reg_layer_2_w23_1), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w24_reg[0] (.CLK(i_clk), .D(n227), .Q(reg_layer_2_w24_0), .Q_N(n141), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w24_reg[1] (.CLK(i_clk), .D(n228), .Q(reg_layer_2_w24_1), .Q_N(n143), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w24_reg[2] (.CLK(i_clk), .D(n229), .Q(reg_layer_2_w24_2), .Q_N(n145), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w25_reg[0] (.CLK(i_clk), .D(n225), .Q(reg_layer_2_w25_0), .Q_N(n137), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w25_reg[1] (.CLK(i_clk), .D(n226), .Q(reg_layer_2_w25_1), .Q_N(n139), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w26_reg[0] (.CLK(i_clk), .D(n222), .Q(reg_layer_2_w26_0), .Q_N(n131), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w26_reg[1] (.CLK(i_clk), .D(n223), .Q(reg_layer_2_w26_1), .Q_N(n133), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w26_reg[2] (.CLK(i_clk), .D(n224), .Q(reg_layer_2_w26_2), .Q_N(n135), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w27_reg[0] (.CLK(i_clk), .D(n220), .Q(reg_layer_2_w27_0), .Q_N(n127), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w27_reg[1] (.CLK(i_clk), .D(n221), .Q(reg_layer_2_w27_1), .Q_N(n129), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w29_reg[0] (.CLK(i_clk), .D(n295), .Q(reg_layer_2_w29_0), .Q_N(n56), .RESET_B(i_rst));
sg13g2_dfrbp_2 \reg_layer_2_w29_reg[1] (.CLK(i_clk), .D(n296), .Q(reg_layer_2_w29_1), .Q_N(n58), .RESET_B(i_rst));
sg13g2_dfrbp_1 \reg_layer_2_w29_reg[2] (.CLK(i_clk), .D(n297), .Q(reg_layer_2_w29_2), .RESET_B(i_rst));
sg13g2_dfrbp_2 reg_layer_2_w1_reg (.CLK(i_clk), .D(n290), .Q(A_1), .Q_N(n47), .RESET_B(i_rst));
sg13g2_dfrbp_2 reg_layer_2_w28_reg (.CLK(i_clk), .D(n219), .Q(layer_4_w28_1), .Q_N(n125), .RESET_B(i_rst));
sg13g2_dfrbp_2 reg_layer_2_w30_reg (.CLK(i_clk), .D(n294), .Q(layer_3_w30_1), .Q_N(n54), .RESET_B(i_rst));
sg13g2_dfrbp_1 reg_layer_2_w31_reg (.CLK(i_clk), .D(n293), .Q(A_31), .RESET_B(i_rst));
sg13g2_dfrbp_1 stage_0_ready_reg (.CLK(i_clk), .D(i_start), .Q(stage_0_ready), .Q_N(n344), .RESET_B(i_rst));
sg13g2_dfrbp_1 stage_1_ready_reg (.CLK(i_clk), .D(stage_0_ready), .Q(o_ready), .RESET_B(i_rst));
sg13g2_o21ai_1 U3 (.A1(stage_0_ready), .A2(n164), .B1(n165), .Y(n239));
sg13g2_nand2_2 U4 (.A(layer_2_w20_2), .B(stage_0_ready), .Y(n165));
sg13g2_o21ai_1 U5 (.A1(n11), .A2(stage_0_ready), .B1(n12), .Y(n272));
sg13g2_nand2_2 U6 (.A(layer_2_w10_1), .B(stage_0_ready), .Y(n12));
sg13g2_nand2_2 U7 (.A(layer_2_w11_1), .B(stage_0_ready), .Y(n4));
sg13g2_inv_2 U9 (.A(n201), .Y(n205));
sg13g2_nand2_2 U10 (.A(layer_2_w11_2), .B(stage_0_ready), .Y(n6));
sg13g2_nand2_2 U11 (.A(layer_2_w8_0), .B(stage_0_ready), .Y(n18));
sg13g2_o21ai_1 U12 (.A1(stage_0_ready), .A2(n9), .B1(n10), .Y(n271));
sg13g2_nand2_2 U13 (.A(layer_1_w11_3), .B(stage_0_ready), .Y(n8));
sg13g2_nand2_2 U15 (.A(layer_2_w10_0), .B(stage_0_ready), .Y(n10));
sg13g2_nand2_2 U16 (.A(layer_2_w25_0), .B(stage_0_ready), .Y(n138));
sg13g2_nand2_2 U18 (.A(layer_2_w23_0), .B(stage_0_ready), .Y(n148));
sg13g2_o21ai_1 U19 (.A1(n211), .A2(stage_0_ready), .B1(n212), .Y(n263));
sg13g2_o21ai_1 U21 (.A1(n125), .A2(stage_0_ready), .B1(n126), .Y(n219));
sg13g2_nand2_2 U22 (.A(n15), .B(reg_layer_2_w14_2), .Y(n19));
sg13g2_o21ai_1 U24 (.A1(n172), .A2(stage_0_ready), .B1(n173), .Y(n243));
sg13g2_o21ai_1 U25 (.A1(n7), .A2(stage_0_ready), .B1(n8), .Y(n270));
sg13g2_o21ai_1 U26 (.A1(n129), .A2(stage_0_ready), .B1(n130), .Y(n221));
sg13g2_o21ai_1 U27 (.A1(n145), .A2(stage_0_ready), .B1(n146), .Y(n229));
sg13g2_o21ai_1 U28 (.A1(n39), .A2(stage_0_ready), .B1(n40), .Y(n286));
sg13g2_o21ai_1 U30 (.A1(n41), .A2(stage_0_ready), .B1(n42), .Y(n287));
sg13g2_nand2_2 U31 (.A(n20), .B(reg_layer_2_w12_1), .Y(n188));
sg13g2_o21ai_1 U32 (.A1(n143), .A2(stage_0_ready), .B1(n144), .Y(n228));
sg13g2_nand2_2 U33 (.A(n338), .B(reg_layer_2_w9_1), .Y(n333));
sg13g2_nand2_2 U34 (.A(n344), .B(reg_layer_2_w11_0), .Y(n332));
sg13g2_o21ai_1 U36 (.A1(n192), .A2(stage_0_ready), .B1(n193), .Y(n253));
sg13g2_nand2_2 U37 (.A(layer_1_w7_3), .B(stage_0_ready), .Y(n24));
sg13g2_o21ai_1 U39 (.A1(n199), .A2(stage_0_ready), .B1(n200), .Y(n257));
sg13g2_nand2_2 U40 (.A(layer_1_w6_0), .B(stage_0_ready), .Y(n26));
sg13g2_o21ai_1 U42 (.A1(n127), .A2(stage_0_ready), .B1(n128), .Y(n220));
sg13g2_nand2_2 U43 (.A(layer_1_w6_1), .B(stage_0_ready), .Y(n28));
sg13g2_o21ai_1 U45 (.A1(n131), .A2(stage_0_ready), .B1(n132), .Y(n222));
sg13g2_nand2_2 U46 (.A(layer_1_w5_0), .B(stage_0_ready), .Y(n30));
sg13g2_o21ai_1 U48 (.A1(n166), .A2(stage_0_ready), .B1(n167), .Y(n240));
sg13g2_nand2_2 U49 (.A(layer_1_w5_1), .B(stage_0_ready), .Y(n32));
sg13g2_o21ai_1 U51 (.A1(n29), .A2(stage_0_ready), .B1(n30), .Y(n281));
sg13g2_nand2_2 U52 (.A(\layer_1_w4[0]), .B(stage_0_ready), .Y(n34));
sg13g2_o21ai_1 U54 (.A1(n43), .A2(stage_0_ready), .B1(n44), .Y(n288));
sg13g2_nand2_2 U55 (.A(negation_2), .B(stage_0_ready), .Y(n36));
sg13g2_o21ai_1 U57 (.A1(n207), .A2(stage_0_ready), .B1(n208), .Y(n261));
sg13g2_nand2_2 U58 (.A(layer_1_w3_0), .B(stage_0_ready), .Y(n38));
sg13g2_nand2_2 U60 (.A(n338), .B(reg_layer_2_w15_0), .Y(n339));
sg13g2_nand2_2 U61 (.A(layer_1_w3_1), .B(stage_0_ready), .Y(n40));
sg13g2_o21ai_1 U63 (.A1(n160), .A2(stage_0_ready), .B1(n161), .Y(n237));
sg13g2_nand2_2 U64 (.A(layer_1_w2_0), .B(stage_0_ready), .Y(n42));
sg13g2_nand2_2 U66 (.A(n344), .B(reg_layer_2_w14_0), .Y(n345));
sg13g2_nand2_2 U67 (.A(layer_1_w2_1), .B(stage_0_ready), .Y(n44));
sg13g2_o21ai_1 U69 (.A1(n213), .A2(stage_0_ready), .B1(n214), .Y(n264));
sg13g2_nand2_2 U70 (.A(negation_1), .B(stage_0_ready), .Y(n46));
sg13g2_o21ai_1 U72 (.A1(n141), .A2(stage_0_ready), .B1(n142), .Y(n227));
sg13g2_nand2_2 U73 (.A(layer_1_w1), .B(stage_0_ready), .Y(n48));
sg13g2_o21ai_1 U75 (.A1(n157), .A2(stage_0_ready), .B1(n158), .Y(n235));
sg13g2_nand2_2 U76 (.A(\layer_1_w0[0]), .B(stage_0_ready), .Y(n50));
sg13g2_o21ai_1 U78 (.A1(n135), .A2(stage_0_ready), .B1(n136), .Y(n224));
sg13g2_nand2_2 U79 (.A(negation_0), .B(stage_0_ready), .Y(n52));
sg13g2_inv_2 U81 (.A(n53), .Y(n293));
sg13g2_nor2_2 U82 (.A(A_31), .B(stage_0_ready), .Y(n53));
sg13g2_o21ai_1 U83 (.A1(n139), .A2(stage_0_ready), .B1(n140), .Y(n226));
sg13g2_nand2_2 U84 (.A(layer_1_w30), .B(stage_0_ready), .Y(n55));
sg13g2_nand2_2 U86 (.A(n15), .B(reg_layer_2_w19_0), .Y(n195));
sg13g2_nand2_2 U87 (.A(\layer_2_w29[0]), .B(stage_0_ready), .Y(n57));
sg13g2_nand2_2 U89 (.A(n20), .B(reg_layer_2_w18_0), .Y(n149));
sg13g2_nand2_2 U90 (.A(\layer_1_w29[0]), .B(stage_0_ready), .Y(n59));
sg13g2_inv_2 U92 (.A(n60), .Y(n297));
sg13g2_nor2_2 U93 (.A(reg_layer_2_w29_2), .B(stage_0_ready), .Y(n60));
sg13g2_o21ai_1 U94 (.A1(i_start), .A2(n61), .B1(n62), .Y(n298));
sg13g2_nand2_2 U95 (.A(i_start), .B(\i_mr[0]), .Y(n62));
sg13g2_o21ai_1 U97 (.A1(i_start), .A2(n63), .B1(n64), .Y(n299));
sg13g2_nand2_2 U98 (.A(\i_mr[1]), .B(i_start), .Y(n64));
sg13g2_o21ai_1 U100 (.A1(i_start), .A2(n65), .B1(n66), .Y(n300));
sg13g2_nand2_2 U101 (.A(\i_mr[2]), .B(i_start), .Y(n66));
sg13g2_o21ai_1 U103 (.A1(i_start), .A2(n67), .B1(n68), .Y(n301));
sg13g2_nand2_2 U104 (.A(\i_mr[3]), .B(i_start), .Y(n68));
sg13g2_o21ai_1 U106 (.A1(i_start), .A2(n69), .B1(n70), .Y(n302));
sg13g2_nand2_2 U107 (.A(\i_mr[4]), .B(i_start), .Y(n70));
sg13g2_o21ai_1 U109 (.A1(i_start), .A2(n71), .B1(n72), .Y(n303));
sg13g2_nand2_2 U110 (.A(\i_mr[5]), .B(i_start), .Y(n72));
sg13g2_o21ai_1 U112 (.A1(i_start), .A2(n73), .B1(n74), .Y(n304));
sg13g2_nand2_2 U113 (.A(\i_mr[6]), .B(i_start), .Y(n74));
sg13g2_o21ai_1 U115 (.A1(i_start), .A2(n75), .B1(n76), .Y(n305));
sg13g2_nand2_2 U116 (.A(\i_mr[7]), .B(i_start), .Y(n76));
sg13g2_o21ai_1 U118 (.A1(i_start), .A2(n77), .B1(n78), .Y(n306));
sg13g2_nand2_2 U119 (.A(\i_mr[8]), .B(i_start), .Y(n78));
sg13g2_o21ai_1 U121 (.A1(i_start), .A2(n79), .B1(n80), .Y(n307));
sg13g2_nand2_2 U122 (.A(\i_mr[9]), .B(i_start), .Y(n80));
sg13g2_o21ai_1 U124 (.A1(i_start), .A2(n81), .B1(n82), .Y(n308));
sg13g2_nand2_2 U125 (.A(\i_mr[10]), .B(i_start), .Y(n82));
sg13g2_o21ai_1 U127 (.A1(i_start), .A2(n83), .B1(n84), .Y(n309));
sg13g2_nand2_2 U128 (.A(\i_mr[11]), .B(i_start), .Y(n84));
sg13g2_o21ai_1 U130 (.A1(i_start), .A2(n85), .B1(n86), .Y(n310));
sg13g2_nand2_2 U131 (.A(\i_mr[12]), .B(i_start), .Y(n86));
sg13g2_o21ai_1 U133 (.A1(i_start), .A2(n87), .B1(n88), .Y(n311));
sg13g2_nand2_2 U134 (.A(\i_mr[13]), .B(i_start), .Y(n88));
sg13g2_o21ai_1 U136 (.A1(i_start), .A2(n89), .B1(n90), .Y(n312));
sg13g2_nand2_2 U137 (.A(\i_mr[14]), .B(i_start), .Y(n90));
sg13g2_o21ai_1 U139 (.A1(i_start), .A2(n91), .B1(n92), .Y(n313));
sg13g2_nand2_2 U140 (.A(\i_mr[15]), .B(i_start), .Y(n92));
sg13g2_o21ai_1 U142 (.A1(i_start), .A2(n93), .B1(n94), .Y(n314));
sg13g2_nand2_2 U143 (.A(\i_md[0]), .B(i_start), .Y(n94));
sg13g2_o21ai_1 U145 (.A1(i_start), .A2(n95), .B1(n96), .Y(n315));
sg13g2_nand2_2 U146 (.A(\i_md[1]), .B(i_start), .Y(n96));
sg13g2_o21ai_1 U148 (.A1(i_start), .A2(n97), .B1(n98), .Y(n316));
sg13g2_nand2_2 U149 (.A(\i_md[2]), .B(i_start), .Y(n98));
sg13g2_o21ai_1 U151 (.A1(i_start), .A2(n99), .B1(n100), .Y(n317));
sg13g2_nand2_2 U152 (.A(\i_md[3]), .B(i_start), .Y(n100));
sg13g2_o21ai_1 U154 (.A1(i_start), .A2(n101), .B1(n102), .Y(n318));
sg13g2_nand2_2 U155 (.A(\i_md[4]), .B(i_start), .Y(n102));
sg13g2_o21ai_1 U157 (.A1(i_start), .A2(n103), .B1(n104), .Y(n319));
sg13g2_nand2_2 U158 (.A(\i_md[5]), .B(i_start), .Y(n104));
sg13g2_o21ai_1 U160 (.A1(i_start), .A2(n105), .B1(n106), .Y(n320));
sg13g2_nand2_2 U161 (.A(\i_md[6]), .B(i_start), .Y(n106));
sg13g2_o21ai_1 U163 (.A1(i_start), .A2(n107), .B1(n108), .Y(n321));
sg13g2_nand2_2 U164 (.A(\i_md[7]), .B(i_start), .Y(n108));
sg13g2_o21ai_1 U166 (.A1(i_start), .A2(n109), .B1(n110), .Y(n322));
sg13g2_nand2_2 U167 (.A(\i_md[8]), .B(i_start), .Y(n110));
sg13g2_o21ai_1 U169 (.A1(i_start), .A2(n111), .B1(n112), .Y(n323));
sg13g2_nand2_2 U170 (.A(\i_md[9]), .B(i_start), .Y(n112));
sg13g2_o21ai_1 U172 (.A1(i_start), .A2(n113), .B1(n114), .Y(n324));
sg13g2_nand2_2 U173 (.A(\i_md[10]), .B(i_start), .Y(n114));
sg13g2_o21ai_1 U175 (.A1(i_start), .A2(n115), .B1(n116), .Y(n325));
sg13g2_nand2_2 U176 (.A(\i_md[11]), .B(i_start), .Y(n116));
sg13g2_o21ai_1 U178 (.A1(i_start), .A2(n117), .B1(n118), .Y(n326));
sg13g2_nand2_2 U179 (.A(\i_md[12]), .B(i_start), .Y(n118));
sg13g2_o21ai_1 U181 (.A1(i_start), .A2(n119), .B1(n120), .Y(n327));
sg13g2_nand2_2 U182 (.A(\i_md[13]), .B(i_start), .Y(n120));
sg13g2_o21ai_1 U184 (.A1(i_start), .A2(n121), .B1(n122), .Y(n328));
sg13g2_nand2_2 U185 (.A(\i_md[14]), .B(i_start), .Y(n122));
sg13g2_o21ai_1 U187 (.A1(i_start), .A2(n123), .B1(n124), .Y(n329));
sg13g2_nand2_2 U188 (.A(\i_md[15]), .B(i_start), .Y(n124));
sg13g2_o21ai_1 U190 (.A1(n184), .A2(stage_0_ready), .B1(n185), .Y(n249));
sg13g2_nand2_2 U191 (.A(n334), .B(reg_layer_2_w16_0), .Y(n335));
sg13g2_o21ai_1 U193 (.A1(n25), .A2(stage_0_ready), .B1(n26), .Y(n279));
sg13g2_nand2_2 U194 (.A(layer_1_w27_0), .B(stage_0_ready), .Y(n128));
sg13g2_o21ai_1 U196 (.A1(n33), .A2(stage_0_ready), .B1(n34), .Y(n283));
sg13g2_nand2_2 U197 (.A(layer_1_w27_1), .B(stage_0_ready), .Y(n130));
sg13g2_o21ai_1 U199 (.A1(n49), .A2(stage_0_ready), .B1(n50), .Y(n291));
sg13g2_nand2_2 U200 (.A(\layer_2_w26[0]), .B(stage_0_ready), .Y(n132));
sg13g2_o21ai_1 U202 (.A1(n54), .A2(stage_0_ready), .B1(n55), .Y(n294));
sg13g2_nand2_2 U203 (.A(layer_1_w26_0), .B(stage_0_ready), .Y(n134));
sg13g2_o21ai_1 U205 (.A1(n56), .A2(stage_0_ready), .B1(n57), .Y(n295));
sg13g2_nand2_2 U206 (.A(layer_1_w26_1), .B(stage_0_ready), .Y(n136));
sg13g2_o21ai_1 U208 (.A1(n17), .A2(stage_0_ready), .B1(n18), .Y(n275));
sg13g2_o21ai_1 U209 (.A1(n209), .A2(stage_0_ready), .B1(n210), .Y(n262));
sg13g2_o21ai_1 U211 (.A1(n137), .A2(stage_0_ready), .B1(n138), .Y(n225));
sg13g2_o21ai_1 U212 (.A1(n13), .A2(stage_0_ready), .B1(n14), .Y(n273));
sg13g2_o21ai_1 U214 (.A1(n133), .A2(stage_0_ready), .B1(n134), .Y(n223));
sg13g2_o21ai_1 U215 (.A1(n155), .A2(stage_0_ready), .B1(n156), .Y(n234));
sg13g2_o21ai_1 U217 (.A1(n162), .A2(stage_0_ready), .B1(n163), .Y(n238));
sg13g2_o21ai_1 U218 (.A1(n170), .A2(stage_0_ready), .B1(n171), .Y(n242));
sg13g2_o21ai_1 U220 (.A1(n176), .A2(stage_0_ready), .B1(n177), .Y(n245));
sg13g2_nand2_2 U221 (.A(layer_1_w24_3), .B(stage_0_ready), .Y(n146));
sg13g2_o21ai_1 U223 (.A1(n180), .A2(stage_0_ready), .B1(n181), .Y(n247));
sg13g2_o21ai_1 U224 (.A1(n186), .A2(stage_0_ready), .B1(n187), .Y(n250));
sg13g2_o21ai_1 U226 (.A1(n190), .A2(stage_0_ready), .B1(n191), .Y(n252));
sg13g2_o21ai_1 U227 (.A1(n197), .A2(stage_0_ready), .B1(n198), .Y(n256));
sg13g2_o21ai_1 U228 (.A1(n203), .A2(stage_0_ready), .B1(n204), .Y(n259));
sg13g2_o21ai_1 U229 (.A1(stage_0_ready), .A2(n151), .B1(n152), .Y(n232));
sg13g2_nand2_2 U230 (.A(layer_2_w22_0), .B(stage_0_ready), .Y(n152));
sg13g2_o21ai_1 U232 (.A1(n217), .A2(stage_0_ready), .B1(n218), .Y(n266));
sg13g2_o21ai_1 U233 (.A1(n3), .A2(stage_0_ready), .B1(n4), .Y(n268));
sg13g2_o21ai_1 U234 (.A1(n23), .A2(stage_0_ready), .B1(n24), .Y(n278));
sg13g2_o21ai_1 U235 (.A1(n27), .A2(stage_0_ready), .B1(n28), .Y(n280));
sg13g2_nand2_2 U236 (.A(layer_2_w21_0), .B(stage_0_ready), .Y(n156));
sg13g2_o21ai_1 U238 (.A1(n31), .A2(stage_0_ready), .B1(n32), .Y(n282));
sg13g2_o21ai_1 U239 (.A1(n35), .A2(stage_0_ready), .B1(n36), .Y(n284));
sg13g2_inv_2 U241 (.A(n159), .Y(n236));
sg13g2_nor2_2 U242 (.A(reg_layer_2_w21_2), .B(stage_0_ready), .Y(n159));
sg13g2_o21ai_1 U243 (.A1(n37), .A2(stage_0_ready), .B1(n38), .Y(n285));
sg13g2_o21ai_1 U244 (.A1(n45), .A2(stage_0_ready), .B1(n46), .Y(n289));
sg13g2_o21ai_1 U246 (.A1(n47), .A2(stage_0_ready), .B1(n48), .Y(n290));
sg13g2_nand2_2 U247 (.A(layer_2_w20_1), .B(stage_0_ready), .Y(n163));
sg13g2_o21ai_1 U249 (.A1(n51), .A2(stage_0_ready), .B1(n52), .Y(n292));
sg13g2_o21ai_1 U250 (.A1(n58), .A2(stage_0_ready), .B1(n59), .Y(n296));
sg13g2_nand2_2 U252 (.A(layer_2_w13_0), .B(stage_0_ready), .Y(n208));
sg13g2_nand2_2 U253 (.A(layer_1_w20_3), .B(stage_0_ready), .Y(n167));
sg13g2_nand2_2 U255 (.A(layer_2_w25_1), .B(stage_0_ready), .Y(n140));
sg13g2_nand2_2 U256 (.A(layer_2_w14_2), .B(stage_0_ready), .Y(n206));
sg13g2_nand2_2 U257 (.A(layer_2_w19_2), .B(stage_0_ready), .Y(n173));
sg13g2_nand2_2 U258 (.A(n154), .B(n1), .Y(n233));
sg13g2_nand2_2 U259 (.A(layer_2_w19_1), .B(stage_0_ready), .Y(n171));
sg13g2_nand2_2 U261 (.A(layer_2_w22_1), .B(stage_0_ready), .Y(n154));
sg13g2_nand2_2 U262 (.A(layer_2_w28), .B(stage_0_ready), .Y(n126));
sg13g2_nand2_2 U264 (.A(layer_2_w20_0), .B(stage_0_ready), .Y(n161));
sg13g2_nand2_2 U265 (.A(n189), .B(n335), .Y(n251));
sg13g2_nand2_2 U266 (.A(layer_2_w9_0), .B(stage_0_ready), .Y(n14));
sg13g2_nand2_2 U267 (.A(layer_2_w14_0), .B(stage_0_ready), .Y(n202));
sg13g2_nand2_2 U268 (.A(layer_2_w18_1), .B(stage_0_ready), .Y(n177));
sg13g2_o21ai_1 U270 (.A1(stage_0_ready), .A2(n178), .B1(n179), .Y(n246));
sg13g2_nand2_2 U271 (.A(layer_2_w18_2), .B(stage_0_ready), .Y(n179));
sg13g2_nand2_2 U273 (.A(n175), .B(n149), .Y(n244));
sg13g2_nand2_2 U274 (.A(layer_1_w18_5), .B(stage_0_ready), .Y(n181));
sg13g2_nand2_2 U276 (.A(layer_2_w15_2), .B(stage_0_ready), .Y(n200));
sg13g2_nand2_2 U277 (.A(layer_2_w12_0), .B(stage_0_ready), .Y(n214));
sg13g2_nand2_2 U279 (.A(n183), .B(n168), .Y(n248));
sg13g2_nand2_2 U280 (.A(layer_2_w17_1), .B(stage_0_ready), .Y(n185));
sg13g2_inv_2 U282 (.A(layer_0_w14_5), .Y(n201));
sg13g2_nand2_2 U283 (.A(n2), .B(n332), .Y(n267));
sg13g2_nand2_2 U285 (.A(layer_2_w11_0), .B(stage_0_ready), .Y(n2));
sg13g2_nand2_2 U286 (.A(layer_2_w9_1), .B(stage_0_ready), .Y(n16));
sg13g2_nand2_2 U287 (.A(layer_2_w24_1), .B(stage_0_ready), .Y(n144));
sg13g2_nand2_2 U288 (.A(reg_layer_2_w22_1), .B(n334), .Y(n1));
sg13g2_nand2_2 U289 (.A(layer_2_w16_1), .B(stage_0_ready), .Y(n191));
sg13g2_mux2_1 U291 (.A0(reg_layer_2_w8_1), .A1(layer_2_w8_1), .S(stage_0_ready), .X(n276));
sg13g2_inv_2 U294 (.A(n194), .Y(n254));
sg13g2_nor2_2 U295 (.A(reg_layer_2_w16_3), .B(stage_0_ready), .Y(n194));
sg13g2_o21ai_1 U296 (.A1(n147), .A2(stage_0_ready), .B1(n148), .Y(n230));
sg13g2_nand2_2 U297 (.A(layer_2_w16_2), .B(stage_0_ready), .Y(n193));
sg13g2_nand2_2 U298 (.A(layer_2_w24_0), .B(stage_0_ready), .Y(n142));
sg13g2_nand2_2 U299 (.A(n202), .B(n345), .Y(n258));
sg13g2_nand2_2 U300 (.A(layer_2_w15_1), .B(stage_0_ready), .Y(n198));
sg13g2_nand2_2 U302 (.A(layer_2_w21_1), .B(stage_0_ready), .Y(n158));
sg13g2_nand2_2 U303 (.A(n169), .B(n195), .Y(n241));
sg13g2_nand2_2 U305 (.A(\layer_2_w7[0]), .B(stage_0_ready), .Y(n22));
sg13g2_nand2_2 U306 (.A(layer_2_w17_2), .B(stage_0_ready), .Y(n187));
sg13g2_nand2_2 U307 (.A(layer_2_w13_1), .B(stage_0_ready), .Y(n210));
sg13g2_nand2_2 U308 (.A(n206), .B(n19), .Y(n260));
sg13g2_nand2_2 U309 (.A(layer_2_w14_1), .B(stage_0_ready), .Y(n204));
sg13g2_inv_2 U311 (.A(stage_0_ready), .Y(n15));
sg13g2_inv_2 U312 (.A(stage_0_ready), .Y(n20));
sg13g2_nand2_2 U313 (.A(n20), .B(n153), .Y(n168));
sg13g2_inv_2 U314 (.A(n182), .Y(n153));
sg13g2_inv_2 U315 (.A(n215), .Y(n330));
sg13g2_nand2_2 U317 (.A(n334), .B(reg_layer_2_w23_1), .Y(n174));
sg13g2_nand2_2 U318 (.A(n174), .B(n150), .Y(n231));
sg13g2_nand2_2 U320 (.A(layer_2_w23_1), .B(stage_0_ready), .Y(n150));
sg13g2_nand2_2 U321 (.A(layer_1_w13_5), .B(stage_0_ready), .Y(n212));
sg13g2_nand2_2 U323 (.A(n216), .B(n188), .Y(n265));
sg13g2_nand2_2 U324 (.A(n16), .B(n333), .Y(n274));
sg13g2_inv_2 U326 (.A(negation_6), .Y(n215));
sg13g2_inv_2 U327 (.A(n340), .Y(n341));
sg13g2_nand2_2 U328 (.A(n15), .B(reg_layer_2_w11_2), .Y(n331));
sg13g2_nand2_2 U329 (.A(n6), .B(n331), .Y(n269));
sg13g2_nand2_2 U330 (.A(layer_1_w12_3), .B(stage_0_ready), .Y(n218));
sg13g2_nand2_2 U332 (.A(layer_2_w12_1), .B(stage_0_ready), .Y(n216));
sg13g2_o21ai_1 U333 (.A1(stage_0_ready), .A2(n21), .B1(n22), .Y(n277));
sg13g2_inv_2 U334 (.A(stage_0_ready), .Y(n334));
sg13g2_inv_2 U335 (.A(negation_3), .Y(n336));
sg13g2_inv_2 U336 (.A(n336), .Y(n337));
sg13g2_nand2_2 U337 (.A(n196), .B(n339), .Y(n255));
sg13g2_inv_2 U338 (.A(stage_0_ready), .Y(n338));
sg13g2_nand2_2 U339 (.A(layer_2_w15_0), .B(stage_0_ready), .Y(n196));
sg13g2_nand2_2 U340 (.A(layer_2_w16_0), .B(stage_0_ready), .Y(n189));
sg13g2_inv_2 U341 (.A(negation_5), .Y(n340));
sg13g2_inv_2 U342 (.A(negation_4), .Y(n342));
sg13g2_inv_2 U343 (.A(n342), .Y(n343));
sg13g2_nand2_2 U345 (.A(layer_2_w18_0), .B(stage_0_ready), .Y(n175));
sg13g2_nand2_2 U346 (.A(layer_2_w17_0), .B(stage_0_ready), .Y(n183));
sg13g2_nand2_2 U347 (.A(layer_2_w19_0), .B(stage_0_ready), .Y(n169));
sg13g2_tiehi U351 (.L_HI(\*Logic1*));
sg13g2_tielo U352 (.L_LO(\*Logic0*));
adder_32bit_1 adder_32bit(.\i_a[0](reg_layer_2_w0_0), .\i_a[1](A_1), .\i_a[2](A_2), .\i_a[3](layer_4_w3_0), .\i_a[4](layer_4_w4_0), .\i_a[5](layer_4_w5_0), .\i_a[6](layer_4_w6_0), .\i_a[7](layer_4_w7_0), .\i_a[8](layer_4_w8_0), .\i_a[9](layer_4_w9_0), .\i_a[10](layer_4_w10_0), .\i_a[11](layer_4_w11_0), .\i_a[12](layer_4_w12_0), .\i_a[13](layer_4_w13_0), .\i_a[14](layer_4_w14_0), .\i_a[15](layer_4_w15_0), .\i_a[16](layer_4_w16_0), .\i_a[17](layer_4_w17_0), .\i_a[18](layer_4_w18_0), .\i_a[19](layer_4_w19_0), .\i_a[20](layer_4_w20_0), .\i_a[21](layer_4_w21_0), .\i_a[22](layer_4_w22_0), .\i_a[23](layer_4_w23_0), .\i_a[24](layer_4_w24_0), .\i_a[25](A_25), .\i_a[26](layer_4_w26_0), .\i_a[27](A_27), .\i_a[28](layer_4_w28_0), .\i_a[29](A_29), .\i_a[30](layer_3_w30_0), .\i_a[31](A_31), .\i_b[0](reg_layer_2_w0_1), .\i_b[1](\*Logic0*), .\i_b[2](\*Logic0*), .\i_b[3](layer_4_w3_1), .\i_b[4](layer_4_w4_1), .\i_b[5](layer_4_w5_1), .\i_b[6](layer_4_w6_1), .\i_b[7](layer_4_w7_1), .\i_b[8](layer_4_w8_1), .\i_b[9](layer_4_w9_1), .\i_b[10](layer_4_w10_1), .\i_b[11](layer_4_w11_1), .\i_b[12](layer_4_w12_1), .\i_b[13](layer_4_w13_1), .\i_b[14](layer_4_w14_1), .\i_b[15](layer_4_w15_1), .\i_b[16](layer_4_w16_1), .\i_b[17](layer_4_w17_1), .\i_b[18](layer_4_w18_1), .\i_b[19](layer_4_w19_1), .\i_b[20](layer_4_w20_1), .\i_b[21](layer_4_w21_1), .\i_b[22](layer_4_w22_1), .\i_b[23](layer_4_w23_1), .\i_b[24](layer_4_w24_1), .\i_b[25](\*Logic0*), .\i_b[26](layer_4_w26_1), .\i_b[27](\*Logic0*), .\i_b[28](layer_4_w28_1), .\i_b[29](\*Logic0*), .\i_b[30](layer_3_w30_1), .\i_b[31](\*Logic0*), .\o_s[0](\o_product[0]), .\o_s[1](\o_product[1]), .\o_s[2](\o_product[2]), .\o_s[3](\o_product[3]), .\o_s[4](\o_product[4]), .\o_s[5](\o_product[5]), .\o_s[6](\o_product[6]), .\o_s[7](\o_product[7]), .\o_s[8](\o_product[8]), .\o_s[9](\o_product[9]), .\o_s[10](\o_product[10]), .\o_s[11](\o_product[11]), .\o_s[12](\o_product[12]), .\o_s[13](\o_product[13]), .\o_s[14](\o_product[14]), .\o_s[15](\o_product[15]), .\o_s[16](\o_product[16]), .\o_s[17](\o_product[17]), .\o_s[18](\o_product[18]), .\o_s[19](\o_product[19]), .\o_s[20](\o_product[20]), .\o_s[21](\o_product[21]), .\o_s[22](\o_product[22]), .\o_s[23](\o_product[23]), .\o_s[24](\o_product[24]), .\o_s[25](\o_product[25]), .\o_s[26](\o_product[26]), .\o_s[27](\o_product[27]), .\o_s[28](\o_product[28]), .\o_s[29](\o_product[29]), .\o_s[30](\o_product[30]), .\o_s[31](\o_product[31]), .i_c(\*Logic0*), .o_c());
booth_array booth_array_0(.\double[0](double_0), .\double[1](double_1), .\double[2](double_2), .\double[3](double_3), .\double[4](double_4), .\double[5](double_5), .\double[6](double_6), .\double[7](double_7), .\multiplier[0](mr_0), .\multiplier[1](mr_1), .\multiplier[2](mr_2), .\multiplier[3](mr_3), .\multiplier[4](mr_4), .\multiplier[5](mr_5), .\multiplier[6](mr_6), .\multiplier[7](mr_7), .\multiplier[8](mr_8), .\multiplier[9](mr_9), .\multiplier[10](mr_10), .\multiplier[11](mr_11), .\multiplier[12](mr_12), .\multiplier[13](mr_13), .\multiplier[14](mr_14), .\multiplier[15](mr_15), .\negation[0](negation_0), .\negation[1](negation_1), .\negation[2](negation_2), .\negation[3](negation_3), .\negation[4](negation_4), .\negation[5](negation_5), .\negation[6](negation_6), .\negation[7](negation_7), .\zero[0](zero_0), .\zero[1](zero_1), .\zero[2](zero_2), .\zero[3](zero_3), .\zero[4](zero_4), .\zero[5](zero_5), .\zero[6](zero_6), .\zero[7](zero_7));
compressor42_0 layer_1_compressor42_0(.A(layer_0_w6_0), .B(layer_0_w6_1), .C(layer_0_w6_2), .carry(layer_1_w7_0), .cin(n337), .cout(layer_1_w7_1), .D(layer_0_w6_3), .S(layer_1_w6_1));
compressor42_1 layer_2_compressor42_7(.A(layer_1_w19_0), .B(layer_1_w19_1), .C(layer_1_w19_2), .carry(layer_2_w20_0), .cin(\*Logic1*), .cout(layer_2_w20_1), .D(layer_1_w19_3), .S(layer_2_w19_2));
compressor42_2 layer_2_compressor42_6(.A(layer_1_w18_0), .B(layer_1_w18_1), .C(layer_1_w18_2), .carry(layer_2_w19_0), .cin(layer_1_w18_4), .cout(layer_2_w19_1), .D(layer_1_w18_3), .S(layer_2_w18_2));
compressor42_3 layer_2_compressor42_5(.A(layer_1_w17_0), .B(layer_1_w17_1), .C(layer_1_w17_2), .carry(layer_2_w18_0), .cin(layer_1_w17_4), .cout(layer_2_w18_1), .D(layer_1_w17_3), .S(layer_2_w17_2));
compressor42_4 layer_2_compressor42_4(.A(layer_1_w16_0), .B(layer_1_w16_1), .C(layer_1_w16_2), .carry(layer_2_w17_0), .cin(layer_1_w16_4), .cout(layer_2_w17_1), .D(layer_1_w16_3), .S(layer_2_w16_2));
compressor42_5 layer_2_compressor42_3(.A(layer_1_w15_0), .B(layer_1_w15_1), .C(layer_1_w15_2), .carry(layer_2_w16_0), .cin(layer_1_w15_4), .cout(layer_2_w16_1), .D(layer_1_w15_3), .S(layer_2_w15_2));
compressor42_6 layer_2_compressor42_2(.A(layer_1_w14_0), .B(layer_1_w14_1), .C(layer_1_w14_2), .carry(layer_2_w15_0), .cin(negation_7), .cout(layer_2_w15_1), .D(layer_1_w14_3), .S(layer_2_w14_2));
compressor42_7 layer_2_compressor42_1(.A(layer_1_w13_0), .B(layer_1_w13_1), .C(layer_1_w13_2), .carry(layer_2_w14_0), .cin(layer_1_w13_4), .cout(layer_2_w14_1), .D(layer_1_w13_3), .S(layer_2_w13_1));
compressor42_8 layer_2_compressor42_0(.A(layer_1_w10_0), .B(layer_1_w10_1), .C(layer_1_w10_2), .carry(layer_2_w11_0), .cin(n341), .cout(layer_2_w11_1), .D(layer_1_w10_3), .S(layer_2_w10_1));
compressor42_9 layer_1_compressor42_16(.A(layer_0_w23_0), .B(layer_0_w23_1), .C(layer_0_w23_2), .carry(layer_1_w24_0), .cin(\*Logic1*), .cout(layer_1_w24_1), .D(layer_0_w23_3), .S(layer_1_w23_2));
compressor42_10 layer_1_compressor42_15(.A(layer_0_w22_0), .B(layer_0_w22_1), .C(layer_0_w22_2), .carry(layer_1_w23_0), .cin(layer_0_w22_4), .cout(layer_1_w23_1), .D(layer_0_w22_3), .S(layer_1_w22_2));
compressor42_11 layer_1_compressor42_14(.A(layer_0_w21_0), .B(layer_0_w21_1), .C(layer_0_w21_2), .carry(layer_1_w22_0), .cin(layer_0_w21_4), .cout(layer_1_w22_1), .D(layer_0_w21_3), .S(layer_1_w21_2));
compressor42_12 layer_1_compressor42_13(.A(layer_0_w20_0), .B(layer_0_w20_1), .C(layer_0_w20_2), .carry(layer_1_w21_0), .cin(layer_0_w20_4), .cout(layer_1_w21_1), .D(layer_0_w20_3), .S(layer_1_w20_2));
compressor42_13 layer_1_compressor42_12(.A(layer_0_w19_0), .B(layer_0_w19_1), .C(layer_0_w19_2), .carry(layer_1_w20_0), .cin(layer_0_w19_4), .cout(layer_1_w20_1), .D(layer_0_w19_3), .S(layer_1_w19_2));
compressor42_14 layer_1_compressor42_11(.A(layer_0_w18_0), .B(layer_0_w18_1), .C(layer_0_w18_2), .carry(layer_1_w19_0), .cin(layer_0_w18_4), .cout(layer_1_w19_1), .D(layer_0_w18_3), .S(layer_1_w18_3));
compressor42_15 layer_1_compressor42_10(.A(layer_0_w17_0), .B(layer_0_w17_1), .C(layer_0_w17_2), .carry(layer_1_w18_0), .cin(layer_0_w17_4), .cout(layer_1_w18_1), .D(layer_0_w17_3), .S(layer_1_w17_3));
compressor42_16 layer_1_compressor42_9(.A(layer_0_w16_0), .B(layer_0_w16_1), .C(layer_0_w16_2), .carry(layer_1_w17_0), .cin(layer_0_w16_4), .cout(layer_1_w17_1), .D(layer_0_w16_3), .S(layer_1_w16_3));
compressor42_17 layer_1_compressor42_8(.A(layer_0_w15_0), .B(layer_0_w15_1), .C(layer_0_w15_2), .carry(layer_1_w16_0), .cin(layer_0_w15_4), .cout(layer_1_w16_1), .D(layer_0_w15_3), .S(layer_1_w15_3));
compressor42_18 layer_1_compressor42_7(.A(layer_0_w14_0), .B(layer_0_w14_1), .C(layer_0_w14_2), .carry(layer_1_w15_0), .cin(layer_0_w14_4), .cout(layer_1_w15_1), .D(layer_0_w14_3), .S(layer_1_w14_2));
compressor42_19 layer_1_compressor42_6(.A(layer_0_w13_0), .B(layer_0_w13_1), .C(layer_0_w13_2), .carry(layer_1_w14_0), .cin(layer_0_w13_4), .cout(layer_1_w14_1), .D(layer_0_w13_3), .S(layer_1_w13_3));
compressor42_20 layer_1_compressor42_5(.A(layer_0_w12_0), .B(layer_0_w12_1), .C(layer_0_w12_2), .carry(layer_1_w13_0), .cin(layer_0_w12_4), .cout(layer_1_w13_1), .D(layer_0_w12_3), .S(layer_1_w12_2));
compressor42_21 layer_1_compressor42_4(.A(layer_0_w11_0), .B(layer_0_w11_1), .C(layer_0_w11_2), .carry(layer_1_w12_0), .cin(layer_0_w11_4), .cout(layer_1_w12_1), .D(layer_0_w11_3), .S(layer_1_w11_2));
compressor42_22 layer_1_compressor42_3(.A(layer_0_w10_0), .B(layer_0_w10_1), .C(layer_0_w10_2), .carry(layer_1_w11_0), .cin(layer_0_w10_4), .cout(layer_1_w11_1), .D(layer_0_w10_3), .S(layer_1_w10_2));
compressor42_23 layer_1_compressor42_2(.A(layer_0_w9_0), .B(layer_0_w9_1), .C(layer_0_w9_2), .carry(layer_1_w10_0), .cin(layer_0_w9_4), .cout(layer_1_w10_1), .D(layer_0_w9_3), .S(layer_1_w9_2));
compressor42_24 layer_1_compressor42_1(.A(layer_0_w8_0), .B(layer_0_w8_1), .C(layer_0_w8_2), .carry(layer_1_w9_0), .cin(layer_0_w8_4), .cout(layer_1_w9_1), .D(layer_0_w8_3), .S(layer_1_w8_1));
full_adder_0 layer_1_full_adder_0(.A(layer_0_w4_0), .B(layer_0_w4_1), .cin(layer_0_w4_2), .cout(layer_1_w5_0), .S(\layer_1_w4[0]));
full_adder_1 layer_4_full_adder_6(.A(\layer_3_w27[0]), .B(reg_layer_2_w27_0), .cin(reg_layer_2_w27_1), .cout(layer_4_w28_0), .S(A_27));
full_adder_2 layer_4_full_adder_5(.A(\layer_3_w25[0]), .B(reg_layer_2_w25_0), .cin(reg_layer_2_w25_1), .cout(layer_4_w26_0), .S(A_25));
full_adder_3 layer_4_full_adder_4(.A(\layer_3_w22[0]), .B(reg_layer_2_w22_0), .cin(reg_layer_2_w22_1), .cout(layer_4_w23_0), .S(layer_4_w22_1));
full_adder_4 layer_4_full_adder_3(.A(layer_3_w20_0), .B(layer_3_w20_1), .cin(reg_layer_2_w20_3), .cout(layer_4_w21_0), .S(layer_4_w20_1));
full_adder_5 layer_4_full_adder_2(.A(layer_3_w18_0), .B(layer_3_w18_1), .cin(reg_layer_2_w18_3), .cout(layer_4_w19_0), .S(layer_4_w18_1));
full_adder_6 layer_4_full_adder_1(.A(layer_3_w16_0), .B(layer_3_w16_1), .cin(reg_layer_2_w16_3), .cout(layer_4_w17_0), .S(layer_4_w16_1));
full_adder_7 layer_4_full_adder_0(.A(reg_layer_2_w2_0), .B(reg_layer_2_w2_1), .cin(reg_layer_2_w2_2), .cout(layer_4_w3_0), .S(A_2));
full_adder_8 layer_3_full_adder_13(.A(reg_layer_2_w29_0), .B(reg_layer_2_w29_1), .cin(reg_layer_2_w29_2), .cout(layer_3_w30_0), .S(A_29));
full_adder_9 layer_3_full_adder_12(.A(reg_layer_2_w26_0), .B(reg_layer_2_w26_1), .cin(reg_layer_2_w26_2), .cout(\layer_3_w27[0]), .S(layer_4_w26_1));
full_adder_10 layer_3_full_adder_11(.A(reg_layer_2_w24_0), .B(reg_layer_2_w24_1), .cin(reg_layer_2_w24_2), .cout(\layer_3_w25[0]), .S(layer_4_w24_1));
full_adder_11 layer_3_full_adder_10(.A(reg_layer_2_w21_0), .B(reg_layer_2_w21_1), .cin(reg_layer_2_w21_2), .cout(\layer_3_w22[0]), .S(layer_3_w21_1));
full_adder_12 layer_3_full_adder_9(.A(reg_layer_2_w20_0), .B(reg_layer_2_w20_1), .cin(reg_layer_2_w20_2), .cout(layer_3_w21_0), .S(layer_3_w20_1));
full_adder_13 layer_3_full_adder_8(.A(reg_layer_2_w19_0), .B(reg_layer_2_w19_1), .cin(reg_layer_2_w19_2), .cout(layer_3_w20_0), .S(layer_3_w19_1));
full_adder_14 layer_3_full_adder_7(.A(reg_layer_2_w18_0), .B(reg_layer_2_w18_1), .cin(reg_layer_2_w18_2), .cout(layer_3_w19_0), .S(layer_3_w18_1));
full_adder_15 layer_3_full_adder_6(.A(reg_layer_2_w17_0), .B(reg_layer_2_w17_1), .cin(reg_layer_2_w17_2), .cout(layer_3_w18_0), .S(layer_3_w17_1));
full_adder_16 layer_3_full_adder_5(.A(reg_layer_2_w16_0), .B(reg_layer_2_w16_1), .cin(reg_layer_2_w16_2), .cout(layer_3_w17_0), .S(layer_3_w16_1));
full_adder_17 layer_3_full_adder_4(.A(reg_layer_2_w15_0), .B(reg_layer_2_w15_1), .cin(reg_layer_2_w15_2), .cout(layer_3_w16_0), .S(layer_3_w15_1));
full_adder_18 layer_3_full_adder_3(.A(reg_layer_2_w14_0), .B(reg_layer_2_w14_1), .cin(reg_layer_2_w14_2), .cout(layer_3_w15_0), .S(layer_3_w14_1));
full_adder_19 layer_3_full_adder_2(.A(reg_layer_2_w13_0), .B(reg_layer_2_w13_1), .cin(reg_layer_2_w13_2), .cout(layer_3_w14_0), .S(layer_3_w13_1));
full_adder_20 layer_3_full_adder_1(.A(reg_layer_2_w12_0), .B(reg_layer_2_w12_1), .cin(reg_layer_2_w12_2), .cout(layer_3_w13_0), .S(layer_3_w12_1));
full_adder_21 layer_3_full_adder_0(.A(reg_layer_2_w11_0), .B(reg_layer_2_w11_1), .cin(reg_layer_2_w11_2), .cout(layer_3_w12_0), .S(\layer_3_w11[0]));
full_adder_22 layer_2_full_adder_11(.A(layer_1_w28_0), .B(layer_1_w28_1), .cin(layer_1_w28_2), .cout(\layer_2_w29[0]), .S(layer_2_w28));
full_adder_23 layer_2_full_adder_10(.A(layer_1_w25_0), .B(layer_1_w25_1), .cin(\*Logic1*), .cout(\layer_2_w26[0]), .S(layer_2_w25_1));
full_adder_24 layer_2_full_adder_9(.A(layer_1_w24_0), .B(layer_1_w24_1), .cin(layer_1_w24_2), .cout(layer_2_w25_0), .S(layer_2_w24_1));
full_adder_25 layer_2_full_adder_8(.A(layer_1_w23_0), .B(layer_1_w23_1), .cin(layer_1_w23_2), .cout(layer_2_w24_0), .S(layer_2_w23_1));
full_adder_26 layer_2_full_adder_7(.A(layer_1_w22_0), .B(layer_1_w22_1), .cin(layer_1_w22_2), .cout(layer_2_w23_0), .S(layer_2_w22_1));
full_adder_27 layer_2_full_adder_6(.A(layer_1_w21_0), .B(layer_1_w21_1), .cin(layer_1_w21_2), .cout(layer_2_w22_0), .S(layer_2_w21_1));
full_adder_28 layer_2_full_adder_5(.A(layer_1_w20_0), .B(layer_1_w20_1), .cin(layer_1_w20_2), .cout(layer_2_w21_0), .S(layer_2_w20_2));
full_adder_29 layer_2_full_adder_4(.A(layer_1_w12_0), .B(layer_1_w12_1), .cin(layer_1_w12_2), .cout(layer_2_w13_0), .S(layer_2_w12_1));
full_adder_30 layer_2_full_adder_3(.A(layer_1_w11_0), .B(layer_1_w11_1), .cin(layer_1_w11_2), .cout(layer_2_w12_0), .S(layer_2_w11_2));
full_adder_31 layer_2_full_adder_2(.A(layer_1_w9_0), .B(layer_1_w9_1), .cin(layer_1_w9_2), .cout(layer_2_w10_0), .S(layer_2_w9_1));
full_adder_32 layer_2_full_adder_1(.A(layer_1_w8_0), .B(layer_1_w8_1), .cin(n343), .cout(layer_2_w9_0), .S(layer_2_w8_1));
full_adder_33 layer_2_full_adder_0(.A(layer_1_w7_0), .B(layer_1_w7_1), .cin(layer_1_w7_2), .cout(layer_2_w8_0), .S(\layer_2_w7[0]));
full_adder_34 layer_1_full_adder_11(.A(layer_0_w27_0), .B(layer_0_w27_1), .cin(\*Logic1*), .cout(layer_1_w28_0), .S(layer_1_w27_1));
full_adder_35 layer_1_full_adder_10(.A(layer_0_w26_0), .B(layer_0_w26_1), .cin(layer_0_w26_2), .cout(layer_1_w27_0), .S(layer_1_w26_1));
full_adder_36 layer_1_full_adder_9(.A(layer_0_w25_0), .B(layer_0_w25_1), .cin(layer_0_w25_2), .cout(layer_1_w26_0), .S(layer_1_w25_1));
full_adder_37 layer_1_full_adder_8(.A(layer_0_w24_0), .B(layer_0_w24_1), .cin(layer_0_w24_2), .cout(layer_1_w25_0), .S(layer_1_w24_2));
full_adder_38 layer_1_full_adder_7(.A(layer_0_w17_5), .B(layer_0_w17_6), .cin(\*Logic1*), .cout(layer_1_w18_2), .S(layer_1_w17_4));
full_adder_39 layer_1_full_adder_6(.A(layer_0_w16_5), .B(layer_0_w16_6), .cin(layer_0_w16_7), .cout(layer_1_w17_2), .S(layer_1_w16_4));
full_adder_40 layer_1_full_adder_5(.A(layer_0_w15_5), .B(layer_0_w15_6), .cin(layer_0_w15_7), .cout(layer_1_w16_2), .S(layer_1_w15_4));
full_adder_41 layer_1_full_adder_4(.A(n205), .B(layer_0_w14_6), .cin(layer_0_w14_7), .cout(layer_1_w15_2), .S(layer_1_w14_3));
full_adder_42 layer_1_full_adder_3(.A(layer_0_w12_5), .B(layer_0_w12_6), .cin(n330), .cout(layer_1_w13_2), .S(layer_1_w12_3));
full_adder_43 layer_1_full_adder_2(.A(layer_0_w7_0), .B(layer_0_w7_1), .cin(layer_0_w7_2), .cout(layer_1_w8_0), .S(layer_1_w7_2));
full_adder_44 layer_1_full_adder_1(.A(layer_0_w5_0), .B(layer_0_w5_1), .cin(layer_0_w5_2), .cout(layer_1_w6_0), .S(layer_1_w5_1));
half_adder_0 layer_4_half_adder_0(.A(reg_layer_2_w3_0), .B(reg_layer_2_w3_1), .carry(layer_4_w4_0), .S(layer_4_w3_1));
half_adder_1 layer_4_half_adder_16(.A(reg_layer_2_w23_0), .B(reg_layer_2_w23_1), .carry(layer_4_w24_0), .S(layer_4_w23_1));
half_adder_2 layer_4_half_adder_15(.A(layer_3_w21_0), .B(layer_3_w21_1), .carry(layer_4_w22_0), .S(layer_4_w21_1));
half_adder_3 layer_4_half_adder_14(.A(layer_3_w19_0), .B(layer_3_w19_1), .carry(layer_4_w20_0), .S(layer_4_w19_1));
half_adder_4 layer_4_half_adder_13(.A(layer_3_w17_0), .B(layer_3_w17_1), .carry(layer_4_w18_0), .S(layer_4_w17_1));
half_adder_5 layer_4_half_adder_12(.A(layer_3_w15_0), .B(layer_3_w15_1), .carry(layer_4_w16_0), .S(layer_4_w15_1));
half_adder_6 layer_4_half_adder_11(.A(layer_3_w14_0), .B(layer_3_w14_1), .carry(layer_4_w15_0), .S(layer_4_w14_1));
half_adder_7 layer_4_half_adder_10(.A(layer_3_w13_0), .B(layer_3_w13_1), .carry(layer_4_w14_0), .S(layer_4_w13_1));
half_adder_8 layer_4_half_adder_9(.A(layer_3_w12_0), .B(layer_3_w12_1), .carry(layer_4_w13_0), .S(layer_4_w12_1));
half_adder_9 layer_4_half_adder_8(.A(\layer_3_w11[0]), .B(reg_layer_2_w11_3), .carry(layer_4_w12_0), .S(layer_4_w11_1));
half_adder_10 layer_4_half_adder_7(.A(reg_layer_2_w10_0), .B(reg_layer_2_w10_1), .carry(layer_4_w11_0), .S(layer_4_w10_1));
half_adder_11 layer_4_half_adder_6(.A(reg_layer_2_w9_0), .B(reg_layer_2_w9_1), .carry(layer_4_w10_0), .S(layer_4_w9_1));
half_adder_12 layer_4_half_adder_5(.A(reg_layer_2_w8_0), .B(reg_layer_2_w8_1), .carry(layer_4_w9_0), .S(layer_4_w8_1));
half_adder_13 layer_4_half_adder_4(.A(reg_layer_2_w7_0), .B(reg_layer_2_w7_1), .carry(layer_4_w8_0), .S(layer_4_w7_1));
half_adder_14 layer_4_half_adder_3(.A(reg_layer_2_w6_0), .B(reg_layer_2_w6_1), .carry(layer_4_w7_0), .S(layer_4_w6_1));
half_adder_15 layer_4_half_adder_2(.A(reg_layer_2_w5_0), .B(reg_layer_2_w5_1), .carry(layer_4_w6_0), .S(layer_4_w5_1));
half_adder_16 layer_4_half_adder_1(.A(reg_layer_2_w4_0), .B(reg_layer_2_w4_1), .carry(layer_4_w5_0), .S(layer_4_w4_1));
partial_product_gen_0 partial_product_gen_0(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](\layer_1_w0[0]), .\pp[1](layer_1_w1), .\pp[2](layer_1_w2_0), .\pp[3](layer_1_w3_0), .\pp[4](layer_0_w4_0), .\pp[5](layer_0_w5_0), .\pp[6](layer_0_w6_0), .\pp[7](layer_0_w7_0), .\pp[8](layer_0_w8_0), .\pp[9](layer_0_w9_0), .\pp[10](layer_0_w10_0), .\pp[11](layer_0_w11_0), .\pp[12](layer_0_w12_0), .\pp[13](layer_0_w13_0), .\pp[14](layer_0_w14_0), .\pp[15](layer_0_w15_0), .\pp[16](layer_0_w16_0), .double(double_0), .negation(negation_0), .zero(zero_0));
partial_product_gen_1 partial_product_gen_7(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_0_w14_7), .\pp[1](layer_0_w15_7), .\pp[2](layer_0_w16_7), .\pp[3](layer_0_w17_6), .\pp[4](layer_1_w18_5), .\pp[5](layer_1_w19_3), .\pp[6](layer_1_w20_3), .\pp[7](layer_0_w21_4), .\pp[8](layer_0_w22_4), .\pp[9](layer_0_w23_3), .\pp[10](layer_1_w24_3), .\pp[11](layer_0_w25_2), .\pp[12](layer_0_w26_2), .\pp[13](layer_0_w27_1), .\pp[14](layer_1_w28_2), .\pp[15](\layer_1_w29[0]), .\pp[16](layer_1_w30), .double(double_7), .negation(negation_7), .zero(zero_7));
partial_product_gen_2 partial_product_gen_6(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_0_w12_6), .\pp[1](layer_1_w13_5), .\pp[2](layer_0_w14_6), .\pp[3](layer_0_w15_6), .\pp[4](layer_0_w16_6), .\pp[5](layer_0_w17_5), .\pp[6](layer_1_w18_4), .\pp[7](layer_0_w19_4), .\pp[8](layer_0_w20_4), .\pp[9](layer_0_w21_3), .\pp[10](layer_0_w22_3), .\pp[11](layer_0_w23_2), .\pp[12](layer_0_w24_2), .\pp[13](layer_0_w25_1), .\pp[14](layer_0_w26_1), .\pp[15](layer_0_w27_0), .\pp[16](layer_1_w28_1), .double(double_6), .negation(n330), .zero(zero_6));
partial_product_gen_3 partial_product_gen_5(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_1_w10_3), .\pp[1](layer_1_w11_3), .\pp[2](layer_0_w12_5), .\pp[3](layer_1_w13_4), .\pp[4](layer_0_w14_5), .\pp[5](layer_0_w15_5), .\pp[6](layer_0_w16_5), .\pp[7](layer_0_w17_4), .\pp[8](layer_0_w18_4), .\pp[9](layer_0_w19_3), .\pp[10](layer_0_w20_3), .\pp[11](layer_0_w21_2), .\pp[12](layer_0_w22_2), .\pp[13](layer_0_w23_1), .\pp[14](layer_0_w24_1), .\pp[15](layer_0_w25_0), .\pp[16](layer_0_w26_0), .double(double_5), .negation(n341), .zero(zero_5));
partial_product_gen_4 partial_product_gen_4(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_0_w8_4), .\pp[1](layer_0_w9_4), .\pp[2](layer_0_w10_4), .\pp[3](layer_0_w11_4), .\pp[4](layer_0_w12_4), .\pp[5](layer_0_w13_4), .\pp[6](layer_0_w14_4), .\pp[7](layer_0_w15_4), .\pp[8](layer_0_w16_4), .\pp[9](layer_0_w17_3), .\pp[10](layer_0_w18_3), .\pp[11](layer_0_w19_2), .\pp[12](layer_0_w20_2), .\pp[13](layer_0_w21_1), .\pp[14](layer_0_w22_1), .\pp[15](layer_0_w23_0), .\pp[16](layer_0_w24_0), .double(double_4), .negation(negation_4), .zero(zero_4));
partial_product_gen_5 partial_product_gen_3(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_0_w6_3), .\pp[1](layer_1_w7_3), .\pp[2](layer_0_w8_3), .\pp[3](layer_0_w9_3), .\pp[4](layer_0_w10_3), .\pp[5](layer_0_w11_3), .\pp[6](layer_0_w12_3), .\pp[7](layer_0_w13_3), .\pp[8](layer_0_w14_3), .\pp[9](layer_0_w15_3), .\pp[10](layer_0_w16_3), .\pp[11](layer_0_w17_2), .\pp[12](layer_0_w18_2), .\pp[13](layer_0_w19_1), .\pp[14](layer_0_w20_1), .\pp[15](layer_0_w21_0), .\pp[16](layer_0_w22_0), .double(double_3), .negation(negation_3), .zero(zero_3));
partial_product_gen_6 partial_product_gen_2(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_0_w4_2), .\pp[1](layer_0_w5_2), .\pp[2](layer_0_w6_2), .\pp[3](layer_0_w7_2), .\pp[4](layer_0_w8_2), .\pp[5](layer_0_w9_2), .\pp[6](layer_0_w10_2), .\pp[7](layer_0_w11_2), .\pp[8](layer_0_w12_2), .\pp[9](layer_0_w13_2), .\pp[10](layer_0_w14_2), .\pp[11](layer_0_w15_2), .\pp[12](layer_0_w16_2), .\pp[13](layer_0_w17_1), .\pp[14](layer_0_w18_1), .\pp[15](layer_0_w19_0), .\pp[16](layer_0_w20_0), .double(double_2), .negation(negation_2), .zero(zero_2));
partial_product_gen_7 partial_product_gen_1(.\md[0](md_0), .\md[1](md_1), .\md[2](md_2), .\md[3](md_3), .\md[4](md_4), .\md[5](md_5), .\md[6](md_6), .\md[7](md_7), .\md[8](md_8), .\md[9](md_9), .\md[10](md_10), .\md[11](md_11), .\md[12](md_12), .\md[13](md_13), .\md[14](md_14), .\md[15](md_15), .\pp[0](layer_1_w2_1), .\pp[1](layer_1_w3_1), .\pp[2](layer_0_w4_1), .\pp[3](layer_0_w5_1), .\pp[4](layer_0_w6_1), .\pp[5](layer_0_w7_1), .\pp[6](layer_0_w8_1), .\pp[7](layer_0_w9_1), .\pp[8](layer_0_w10_1), .\pp[9](layer_0_w11_1), .\pp[10](layer_0_w12_1), .\pp[11](layer_0_w13_1), .\pp[12](layer_0_w14_1), .\pp[13](layer_0_w15_1), .\pp[14](layer_0_w16_1), .\pp[15](layer_0_w17_0), .\pp[16](layer_0_w18_0), .double(double_1), .negation(negation_1), .zero(zero_1));
endmodule

module adder_32bit_1 (\i_a[0], \i_a[1], \i_a[2], \i_a[3], \i_a[4], \i_a[5], \i_a[6], \i_a[7], \i_a[8], \i_a[9], \i_a[10], \i_a[11], \i_a[12], \i_a[13], \i_a[14], \i_a[15], \i_a[16], \i_a[17], \i_a[18], \i_a[19], \i_a[20], \i_a[21], \i_a[22], \i_a[23], \i_a[24], \i_a[25], \i_a[26], \i_a[27], \i_a[28], \i_a[29], \i_a[30], \i_a[31], \i_b[0], \i_b[1], \i_b[2], \i_b[3], \i_b[4], \i_b[5], \i_b[6], \i_b[7], \i_b[8], \i_b[9], \i_b[10], \i_b[11], \i_b[12], \i_b[13], \i_b[14], \i_b[15], \i_b[16], \i_b[17], \i_b[18], \i_b[19], \i_b[20], \i_b[21], \i_b[22], \i_b[23], \i_b[24], \i_b[25], \i_b[26], \i_b[27], \i_b[28], \i_b[29], \i_b[30], \i_b[31], \o_s[0], \o_s[1], \o_s[2], \o_s[3], \o_s[4], \o_s[5], \o_s[6], \o_s[7], \o_s[8], \o_s[9], \o_s[10], \o_s[11], \o_s[12], \o_s[13], \o_s[14], \o_s[15], \o_s[16], \o_s[17], \o_s[18], \o_s[19], \o_s[20], \o_s[21], \o_s[22], \o_s[23], \o_s[24], \o_s[25], \o_s[26], \o_s[27], \o_s[28], \o_s[29], \o_s[30], \o_s[31], i_c, o_c);
input \i_a[0], \i_a[1], \i_a[2], \i_a[3], \i_a[4], \i_a[5], \i_a[6], \i_a[7], \i_a[8], \i_a[9], \i_a[10], \i_a[11], \i_a[12], \i_a[13], \i_a[14], \i_a[15], \i_a[16], \i_a[17], \i_a[18], \i_a[19], \i_a[20], \i_a[21], \i_a[22], \i_a[23], \i_a[24], \i_a[25], \i_a[26], \i_a[27], \i_a[28], \i_a[29], \i_a[30], \i_a[31], \i_b[0], \i_b[1], \i_b[2], \i_b[3], \i_b[4], \i_b[5], \i_b[6], \i_b[7], \i_b[8], \i_b[9], \i_b[10], \i_b[11], \i_b[12], \i_b[13], \i_b[14], \i_b[15], \i_b[16], \i_b[17], \i_b[18], \i_b[19], \i_b[20], \i_b[21], \i_b[22], \i_b[23], \i_b[24], \i_b[25], \i_b[26], \i_b[27], \i_b[28], \i_b[29], \i_b[30], \i_b[31], i_c;
output \o_s[0], \o_s[1], \o_s[2], \o_s[3], \o_s[4], \o_s[5], \o_s[6], \o_s[7], \o_s[8], \o_s[9], \o_s[10], \o_s[11], \o_s[12], \o_s[13], \o_s[14], \o_s[15], \o_s[16], \o_s[17], \o_s[18], \o_s[19], \o_s[20], \o_s[21], \o_s[22], \o_s[23], \o_s[24], \o_s[25], \o_s[26], \o_s[27], \o_s[28], \o_s[29], \o_s[30], \o_s[31], o_c;

sg13g2_inv_2 U1 (.A(n93), .Y(\o_s[9]));
sg13g2_xnor2_1 U2 (.A(P0_9), .B(G4_4), .Y(n93));
sg13g2_inv_2 U3 (.A(n92), .Y(\o_s[8]));
sg13g2_xnor2_1 U4 (.A(n58), .B(G6_7), .Y(n92));
sg13g2_inv_2 U5 (.A(n91), .Y(\o_s[7]));
sg13g2_xnor2_1 U6 (.A(P0_7), .B(G3_3), .Y(n91));
sg13g2_inv_2 U7 (.A(n90), .Y(\o_s[6]));
sg13g2_xnor2_1 U8 (.A(P0_6), .B(G6_5), .Y(n90));
sg13g2_inv_2 U9 (.A(n89), .Y(\o_s[5]));
sg13g2_xnor2_1 U10 (.A(P0_5), .B(G3_2), .Y(n89));
sg13g2_inv_2 U11 (.A(n88), .Y(\o_s[4]));
sg13g2_xnor2_1 U12 (.A(P0_4), .B(G6_3), .Y(n88));
sg13g2_inv_2 U13 (.A(n87), .Y(\o_s[3]));
sg13g2_xnor2_1 U14 (.A(P0_3), .B(G2_1), .Y(n87));
sg13g2_inv_2 U15 (.A(n77), .Y(\o_s[16]));
sg13g2_buf_2 U16 (.A(G4_7), .X(n8));
sg13g2_xnor2_1 U17 (.A(n9), .B(n14), .Y(n85));
sg13g2_inv_2 U18 (.A(P0_29), .Y(n9));
sg13g2_inv_2 U19 (.A(n86), .Y(\o_s[2]));
sg13g2_xnor2_1 U20 (.A(P0_2), .B(G6_1), .Y(n86));
sg13g2_inv_2 U21 (.A(G5_14), .Y(n14));
sg13g2_xnor2_1 U22 (.A(n18), .B(\G6[29]), .Y(\o_s[30]));
sg13g2_inv_2 U23 (.A(P0_30), .Y(n18));
sg13g2_xnor2_1 U24 (.A(G5_9), .B(P0_19), .Y(n78));
sg13g2_inv_2 U25 (.A(P0_24), .Y(n36));
sg13g2_inv_2 U26 (.A(P0_31), .Y(n55));
sg13g2_nand2_2 U27 (.A(n40), .B(n39), .Y(n82));
sg13g2_nand2_2 U28 (.A(G5_12), .B(P0_25), .Y(n39));
sg13g2_xnor2_1 U29 (.A(G5_8), .B(n67), .Y(\o_s[17]));
sg13g2_inv_2 U30 (.A(n74), .Y(\o_s[12]));
sg13g2_inv_2 U31 (.A(n83), .Y(\o_s[27]));
sg13g2_nand2_2 U32 (.A(n35), .B(n34), .Y(n20));
sg13g2_inv_2 U33 (.A(n20), .Y(\o_s[20]));
sg13g2_nand2_2 U34 (.A(G6_19), .B(n24), .Y(n34));
sg13g2_inv_2 U35 (.A(n27), .Y(n24));
sg13g2_inv_2 U36 (.A(P0_20), .Y(n27));
sg13g2_inv_2 U37 (.A(n80), .Y(\o_s[21]));
sg13g2_xnor2_1 U38 (.A(P0_21), .B(G5_10), .Y(n80));
sg13g2_nand2_2 U39 (.A(n33), .B(n27), .Y(n35));
sg13g2_inv_2 U40 (.A(G6_19), .Y(n33));
sg13g2_inv_2 U41 (.A(n79), .Y(\o_s[1]));
sg13g2_xnor2_1 U42 (.A(P0_1), .B(G1_0), .Y(n79));
sg13g2_xnor2_1 U43 (.A(n36), .B(G6_23), .Y(\o_s[24]));
sg13g2_xnor2_1 U44 (.A(n59), .B(G6_21), .Y(\o_s[22]));
sg13g2_inv_2 U45 (.A(n84), .Y(\o_s[28]));
sg13g2_nand2_2 U46 (.A(n37), .B(n38), .Y(n40));
sg13g2_inv_2 U47 (.A(G5_12), .Y(n37));
sg13g2_inv_2 U48 (.A(P0_25), .Y(n38));
sg13g2_inv_2 U49 (.A(n82), .Y(\o_s[25]));
sg13g2_xnor2_1 U50 (.A(n62), .B(G6_17), .Y(\o_s[18]));
sg13g2_inv_2 U51 (.A(n76), .Y(\o_s[15]));
sg13g2_xnor2_1 U52 (.A(G4_7), .B(n70), .Y(n76));
sg13g2_inv_2 U53 (.A(G0_13), .Y(n42));
sg13g2_inv_2 U54 (.A(n42), .Y(n43));
sg13g2_inv_2 U55 (.A(n75), .Y(\o_s[13]));
sg13g2_xnor2_1 U56 (.A(G4_6), .B(P0_13), .Y(n75));
sg13g2_xnor2_1 U57 (.A(n45), .B(G6_25), .Y(\o_s[26]));
sg13g2_inv_2 U58 (.A(P0_26), .Y(n45));
sg13g2_inv_2 U59 (.A(n73), .Y(\o_s[11]));
sg13g2_xnor2_1 U60 (.A(G4_5), .B(P0_11), .Y(n73));
sg13g2_inv_2 U61 (.A(n72), .Y(\o_s[10]));
sg13g2_xnor2_1 U62 (.A(P0_10), .B(G6_9), .Y(n72));
sg13g2_inv_2 U63 (.A(n71), .Y(\o_s[0]));
sg13g2_xnor2_1 U64 (.A(i_c), .B(P0_0), .Y(n71));
sg13g2_nand2_2 U65 (.A(G5_11), .B(P0_23), .Y(n48));
sg13g2_nand2_2 U66 (.A(n47), .B(n46), .Y(n49));
sg13g2_nand2_2 U67 (.A(n48), .B(n49), .Y(n81));
sg13g2_inv_2 U68 (.A(P0_23), .Y(n46));
sg13g2_inv_2 U69 (.A(G5_11), .Y(n47));
sg13g2_inv_2 U70 (.A(n81), .Y(\o_s[23]));
sg13g2_xnor2_1 U71 (.A(n51), .B(G6_11), .Y(n74));
sg13g2_inv_2 U72 (.A(P0_12), .Y(n50));
sg13g2_inv_2 U73 (.A(n50), .Y(n51));
sg13g2_xnor2_1 U74 (.A(n61), .B(G6_15), .Y(n77));
sg13g2_xnor2_1 U75 (.A(G6_13), .B(n66), .Y(\o_s[14]));
sg13g2_xnor2_1 U76 (.A(n55), .B(G5_15), .Y(\o_s[31]));
sg13g2_xnor2_1 U77 (.A(P0_27), .B(G5_13), .Y(n83));
sg13g2_buf_2 U78 (.A(P2_4), .X(n56));
sg13g2_inv_2 U79 (.A(P0_8), .Y(n57));
sg13g2_inv_2 U80 (.A(n57), .Y(n58));
sg13g2_inv_2 U81 (.A(n85), .Y(\o_s[29]));
sg13g2_inv_2 U82 (.A(P0_22), .Y(n59));
sg13g2_inv_2 U83 (.A(P0_16), .Y(n60));
sg13g2_inv_2 U84 (.A(n60), .Y(n61));
sg13g2_inv_2 U85 (.A(n78), .Y(\o_s[19]));
sg13g2_xnor2_1 U86 (.A(n63), .B(G6_27), .Y(n84));
sg13g2_inv_2 U87 (.A(P0_18), .Y(n62));
sg13g2_inv_2 U88 (.A(n67), .Y(n68));
sg13g2_buf_2 U89 (.A(P0_28), .X(n63));
sg13g2_inv_2 U90 (.A(G0_17), .Y(n64));
sg13g2_inv_2 U91 (.A(n64), .Y(n65));
sg13g2_inv_2 U92 (.A(P0_14), .Y(n66));
sg13g2_inv_2 U93 (.A(P0_17), .Y(n67));
sg13g2_inv_2 U94 (.A(P0_15), .Y(n69));
sg13g2_inv_2 U95 (.A(n69), .Y(n70));
operator_A_1 operator_A_31(.A(\i_a[31]), .B(\i_b[31]), .G(G0_31), .P(P0_31));
operator_A_2 operator_A_30(.A(\i_a[30]), .B(\i_b[30]), .G(G0_30), .P(P0_30));
operator_A_3 operator_A_29(.A(\i_a[29]), .B(\i_b[29]), .G(G0_29), .P(P0_29));
operator_A_4 operator_A_28(.A(\i_a[28]), .B(\i_b[28]), .G(G0_28), .P(P0_28));
operator_A_5 operator_A_27(.A(\i_a[27]), .B(\i_b[27]), .G(G0_27), .P(P0_27));
operator_A_6 operator_A_26(.A(\i_a[26]), .B(\i_b[26]), .G(G0_26), .P(P0_26));
operator_A_7 operator_A_25(.A(\i_a[25]), .B(\i_b[25]), .G(G0_25), .P(P0_25));
operator_A_8 operator_A_24(.A(\i_a[24]), .B(\i_b[24]), .G(G0_24), .P(P0_24));
operator_A_9 operator_A_23(.A(\i_a[23]), .B(\i_b[23]), .G(G0_23), .P(P0_23));
operator_A_10 operator_A_22(.A(\i_a[22]), .B(\i_b[22]), .G(G0_22), .P(P0_22));
operator_A_11 operator_A_21(.A(\i_a[21]), .B(\i_b[21]), .G(G0_21), .P(P0_21));
operator_A_12 operator_A_20(.A(\i_a[20]), .B(\i_b[20]), .G(G0_20), .P(P0_20));
operator_A_13 operator_A_19(.A(\i_a[19]), .B(\i_b[19]), .G(G0_19), .P(P0_19));
operator_A_14 operator_A_18(.A(\i_a[18]), .B(\i_b[18]), .G(G0_18), .P(P0_18));
operator_A_15 operator_A_17(.A(\i_a[17]), .B(\i_b[17]), .G(G0_17), .P(P0_17));
operator_A_16 operator_A_16(.A(\i_a[16]), .B(\i_b[16]), .G(G0_16), .P(P0_16));
operator_A_17 operator_A_15(.A(\i_a[15]), .B(\i_b[15]), .G(G0_15), .P(P0_15));
operator_A_18 operator_A_14(.A(\i_a[14]), .B(\i_b[14]), .G(G0_14), .P(P0_14));
operator_A_19 operator_A_13(.A(\i_a[13]), .B(\i_b[13]), .G(G0_13), .P(P0_13));
operator_A_20 operator_A_12(.A(\i_a[12]), .B(\i_b[12]), .G(G0_12), .P(P0_12));
operator_A_21 operator_A_11(.A(\i_a[11]), .B(\i_b[11]), .G(G0_11), .P(P0_11));
operator_A_22 operator_A_10(.A(\i_a[10]), .B(\i_b[10]), .G(G0_10), .P(P0_10));
operator_A_23 operator_A_9(.A(\i_a[9]), .B(\i_b[9]), .G(G0_9), .P(P0_9));
operator_A_24 operator_A_8(.A(\i_a[8]), .B(\i_b[8]), .G(G0_8), .P(P0_8));
operator_A_25 operator_A_7(.A(\i_a[7]), .B(\i_b[7]), .G(G0_7), .P(P0_7));
operator_A_26 operator_A_6(.A(\i_a[6]), .B(\i_b[6]), .G(G0_6), .P(P0_6));
operator_A_27 operator_A_5(.A(\i_a[5]), .B(\i_b[5]), .G(G0_5), .P(P0_5));
operator_A_28 operator_A_4(.A(\i_a[4]), .B(\i_b[4]), .G(G0_4), .P(P0_4));
operator_A_29 operator_A_3(.A(\i_a[3]), .B(\i_b[3]), .G(G0_3), .P(P0_3));
operator_A_30 operator_A_2(.A(\i_a[2]), .B(\i_b[2]), .G(G0_2), .P(P0_2));
operator_A_31 operator_A_1(.A(\i_a[1]), .B(\i_b[1]), .G(G0_1), .P(P0_1));
operator_A_32 operator_A_0(.A(\i_a[0]), .B(\i_b[0]), .G(G0_0), .P(P0_0));
operator_B_1 operator_B_stage_4_15(.G(G3_15), .G1(G3_11), .Go(G4_15), .P(P3_15), .P1(P3_11), .Po(P4_15));
operator_B_2 operator_B_stage_4_14(.G(G3_14), .G1(G3_10), .Go(G4_14), .P(P3_14), .P1(P3_10), .Po(P4_14));
operator_B_3 operator_B_stage_4_13(.G(G3_13), .G1(G3_9), .Go(G4_13), .P(P3_13), .P1(P3_9), .Po(P4_13));
operator_B_4 operator_B_stage_4_12(.G(G3_12), .G1(G3_8), .Go(G4_12), .P(P3_12), .P1(P3_8), .Po(P4_12));
operator_B_5 operator_B_stage_4_11(.G(G3_11), .G1(G3_7), .Go(G4_11), .P(P3_11), .P1(P3_7), .Po(P4_11));
operator_B_6 operator_B_stage_4_10(.G(G3_10), .G1(G3_6), .Go(G4_10), .P(P3_10), .P1(P3_6), .Po(P4_10));
operator_B_7 operator_B_stage_4_9(.G(G3_9), .G1(G3_5), .Go(G4_9), .P(P3_9), .P1(P3_5), .Po(P4_9));
operator_B_8 operator_B_stage_4_8(.G(G3_8), .G1(G3_4), .Go(G4_8), .P(P3_8), .P1(P3_4), .Po(P4_8));
operator_B_9 operator_B_stage_3_15(.G(G2_15), .G1(G2_13), .Go(G3_15), .P(P2_15), .P1(P2_13), .Po(P3_15));
operator_B_10 operator_B_stage_3_14(.G(G2_14), .G1(G2_12), .Go(G3_14), .P(P2_14), .P1(P2_12), .Po(P3_14));
operator_B_11 operator_B_stage_3_13(.G(G2_13), .G1(G2_11), .Go(G3_13), .P(P2_13), .P1(P2_11), .Po(P3_13));
operator_B_12 operator_B_stage_3_12(.G(G2_12), .G1(G2_10), .Go(G3_12), .P(P2_12), .P1(P2_10), .Po(P3_12));
operator_B_13 operator_B_stage_3_11(.G(G2_11), .G1(G2_9), .Go(G3_11), .P(P2_11), .P1(P2_9), .Po(P3_11));
operator_B_14 operator_B_stage_3_10(.G(G2_10), .G1(G2_8), .Go(G3_10), .P(P2_10), .P1(P2_8), .Po(P3_10));
operator_B_15 operator_B_stage_3_9(.G(G2_9), .G1(G2_7), .Go(G3_9), .P(P2_9), .P1(P2_7), .Po(P3_9));
operator_B_16 operator_B_stage_3_8(.G(G2_8), .G1(G2_6), .Go(G3_8), .P(P2_8), .P1(P2_6), .Po(P3_8));
operator_B_17 operator_B_stage_3_7(.G(G2_7), .G1(G2_5), .Go(G3_7), .P(P2_7), .P1(P2_5), .Po(P3_7));
operator_B_18 operator_B_stage_3_6(.G(G2_6), .G1(G2_4), .Go(G3_6), .P(P2_6), .P1(n56), .Po(P3_6));
operator_B_19 operator_B_stage_3_5(.G(G2_5), .G1(G2_3), .Go(G3_5), .P(P2_5), .P1(P2_3), .Po(P3_5));
operator_B_20 operator_B_stage_3_4(.G(G2_4), .G1(G2_2), .Go(G3_4), .P(P2_4), .P1(P2_2), .Po(P3_4));
operator_B_21 operator_B_stage_2_15(.G(G1_15), .G1(G1_14), .Go(G2_15), .P(P1_15), .P1(P1_14), .Po(P2_15));
operator_B_22 operator_B_stage_2_14(.G(G1_14), .G1(G1_13), .Go(G2_14), .P(P1_14), .P1(P1_13), .Po(P2_14));
operator_B_23 operator_B_stage_2_13(.G(G1_13), .G1(G1_12), .Go(G2_13), .P(P1_13), .P1(P1_12), .Po(P2_13));
operator_B_24 operator_B_stage_2_12(.G(G1_12), .G1(G1_11), .Go(G2_12), .P(P1_12), .P1(P1_11), .Po(P2_12));
operator_B_25 operator_B_stage_2_11(.G(G1_11), .G1(G1_10), .Go(G2_11), .P(P1_11), .P1(P1_10), .Po(P2_11));
operator_B_26 operator_B_stage_2_10(.G(G1_10), .G1(G1_9), .Go(G2_10), .P(P1_10), .P1(P1_9), .Po(P2_10));
operator_B_27 operator_B_stage_2_9(.G(G1_9), .G1(G1_8), .Go(G2_9), .P(P1_9), .P1(P1_8), .Po(P2_9));
operator_B_28 operator_B_stage_2_8(.G(G1_8), .G1(G1_7), .Go(G2_8), .P(P1_8), .P1(P1_7), .Po(P2_8));
operator_B_29 operator_B_stage_2_7(.G(G1_7), .G1(G1_6), .Go(G2_7), .P(P1_7), .P1(P1_6), .Po(P2_7));
operator_B_30 operator_B_stage_2_6(.G(G1_6), .G1(G1_5), .Go(G2_6), .P(P1_6), .P1(P1_5), .Po(P2_6));
operator_B_31 operator_B_stage_2_5(.G(G1_5), .G1(G1_4), .Go(G2_5), .P(P1_5), .P1(P1_4), .Po(P2_5));
operator_B_32 operator_B_stage_2_4(.G(G1_4), .G1(G1_3), .Go(G2_4), .P(P1_4), .P1(P1_3), .Po(P2_4));
operator_B_33 operator_B_stage_2_3(.G(G1_3), .G1(G1_2), .Go(G2_3), .P(P1_3), .P1(P1_2), .Po(P2_3));
operator_B_34 operator_B_stage_2_2(.G(G1_2), .G1(G1_1), .Go(G2_2), .P(P1_2), .P1(P1_1), .Po(P2_2));
operator_B_35 operator_B_stage_1_15(.G(G0_30), .G1(G0_29), .Go(G1_15), .P(P0_30), .P1(P0_29), .Po(P1_15));
operator_B_36 operator_B_stage_1_14(.G(G0_28), .G1(G0_27), .Go(G1_14), .P(n63), .P1(P0_27), .Po(P1_14));
operator_B_37 operator_B_stage_1_13(.G(G0_26), .G1(G0_25), .Go(G1_13), .P(P0_26), .P1(P0_25), .Po(P1_13));
operator_B_38 operator_B_stage_1_12(.G(G0_24), .G1(G0_23), .Go(G1_12), .P(P0_24), .P1(P0_23), .Po(P1_12));
operator_B_39 operator_B_stage_1_11(.G(G0_22), .G1(G0_21), .Go(G1_11), .P(P0_22), .P1(P0_21), .Po(P1_11));
operator_B_40 operator_B_stage_1_10(.G(G0_20), .G1(G0_19), .Go(G1_10), .P(P0_20), .P1(P0_19), .Po(P1_10));
operator_B_41 operator_B_stage_1_9(.G(G0_18), .G1(G0_17), .Go(G1_9), .P(P0_18), .P1(P0_17), .Po(P1_9));
operator_B_42 operator_B_stage_1_8(.G(G0_16), .G1(G0_15), .Go(G1_8), .P(P0_16), .P1(P0_15), .Po(P1_8));
operator_B_43 operator_B_stage_1_7(.G(G0_14), .G1(G0_13), .Go(G1_7), .P(P0_14), .P1(P0_13), .Po(P1_7));
operator_B_44 operator_B_stage_1_6(.G(G0_12), .G1(G0_11), .Go(G1_6), .P(P0_12), .P1(P0_11), .Po(P1_6));
operator_B_45 operator_B_stage_1_5(.G(G0_10), .G1(G0_9), .Go(G1_5), .P(P0_10), .P1(P0_9), .Po(P1_5));
operator_B_46 operator_B_stage_1_4(.G(G0_8), .G1(G0_7), .Go(G1_4), .P(P0_8), .P1(P0_7), .Po(P1_4));
operator_B_47 operator_B_stage_1_3(.G(G0_6), .G1(G0_5), .Go(G1_3), .P(P0_6), .P1(P0_5), .Po(P1_3));
operator_B_48 operator_B_stage_1_2(.G(G0_4), .G1(G0_3), .Go(G1_2), .P(P0_4), .P1(P0_3), .Po(P1_2));
operator_B_49 operator_B_stage_1_1(.G(G0_2), .G1(G0_1), .Go(G1_1), .P(P0_2), .P1(P0_1), .Po(P1_1));
operator_C_1 operator_C_stage_6_15(.G(G0_31), .G1(G5_15), .Go(o_c), .P(P0_31));
operator_C_2 operator_C_stage_6_14(.G(G0_29), .G1(G5_14), .Go(\G6[29]), .P(P0_29));
operator_C_3 operator_C_stage_6_13(.G(G0_27), .G1(G5_13), .Go(G6_27), .P(P0_27));
operator_C_4 operator_C_stage_6_12(.G(G0_25), .G1(G5_12), .Go(G6_25), .P(P0_25));
operator_C_5 operator_C_stage_6_11(.G(G0_23), .G1(G5_11), .Go(G6_23), .P(P0_23));
operator_C_6 operator_C_stage_6_10(.G(G0_21), .G1(G5_10), .Go(G6_21), .P(P0_21));
operator_C_7 operator_C_stage_6_9(.G(G0_19), .G1(G5_9), .Go(G6_19), .P(P0_19));
operator_C_8 operator_C_stage_6_8(.G(n65), .G1(G5_8), .Go(G6_17), .P(n68));
operator_C_9 operator_C_stage_6_7(.G(G0_15), .G1(G4_7), .Go(G6_15), .P(n70));
operator_C_10 operator_C_stage_6_6(.G(n43), .G1(G4_6), .Go(G6_13), .P(P0_13));
operator_C_11 operator_C_stage_6_5(.G(G0_11), .G1(G4_5), .Go(G6_11), .P(P0_11));
operator_C_12 operator_C_stage_6_4(.G(G0_9), .G1(G4_4), .Go(G6_9), .P(P0_9));
operator_C_13 operator_C_stage_6_3(.G(G0_7), .G1(G3_3), .Go(G6_7), .P(P0_7));
operator_C_14 operator_C_stage_6_2(.G(G0_5), .G1(G3_2), .Go(G6_5), .P(P0_5));
operator_C_15 operator_C_stage_6_1(.G(G0_3), .G1(G2_1), .Go(G6_3), .P(P0_3));
operator_C_16 operator_C_stage_6_0(.G(G0_1), .G1(G1_0), .Go(G6_1), .P(P0_1));
operator_C_17 operator_C_stage_5_15(.G(G4_15), .G1(n8), .Go(G5_15), .P(P4_15));
operator_C_18 operator_C_stage_5_14(.G(G4_14), .G1(G4_6), .Go(G5_14), .P(P4_14));
operator_C_19 operator_C_stage_5_13(.G(G4_13), .G1(G4_5), .Go(G5_13), .P(P4_13));
operator_C_20 operator_C_stage_5_12(.G(G4_12), .G1(G4_4), .Go(G5_12), .P(P4_12));
operator_C_21 operator_C_stage_5_11(.G(G4_11), .G1(G3_3), .Go(G5_11), .P(P4_11));
operator_C_22 operator_C_stage_5_10(.G(G4_10), .G1(G3_2), .Go(G5_10), .P(P4_10));
operator_C_23 operator_C_stage_5_9(.G(G4_9), .G1(G2_1), .Go(G5_9), .P(P4_9));
operator_C_24 operator_C_stage_5_8(.G(G4_8), .G1(G1_0), .Go(G5_8), .P(P4_8));
operator_C_25 operator_C_stage_4_7(.G(G3_7), .G1(G3_3), .Go(G4_7), .P(P3_7));
operator_C_26 operator_C_stage_4_6(.G(G3_6), .G1(G3_2), .Go(G4_6), .P(P3_6));
operator_C_27 operator_C_stage_4_5(.G(G3_5), .G1(G2_1), .Go(G4_5), .P(P3_5));
operator_C_28 operator_C_stage_4_4(.G(G3_4), .G1(G1_0), .Go(G4_4), .P(P3_4));
operator_C_29 operator_C_stage_3_3(.G(G2_3), .G1(G2_1), .Go(G3_3), .P(P2_3));
operator_C_30 operator_C_stage_3_2(.G(G2_2), .G1(G1_0), .Go(G3_2), .P(P2_2));
operator_C_31 operator_C_stage_2_1(.G(G1_1), .G1(G1_0), .Go(G2_1), .P(P1_1));
operator_C_32 operator_C_stage_1_0(.G(G0_0), .G1(i_c), .Go(G1_0), .P(P0_0));
endmodule

module operator_A_1 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_2 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_3 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_4 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(B), .Y(n6));
sg13g2_nand2_2 U2 (.A(A), .B(n6), .Y(n3));
sg13g2_inv_2 U3 (.A(n7), .Y(G));
sg13g2_nand2_2 U4 (.A(n1), .B(B), .Y(n4));
sg13g2_nand2_2 U5 (.A(n4), .B(n3), .Y(P));
sg13g2_inv_2 U6 (.A(A), .Y(n1));
sg13g2_nand2_2 U7 (.A(A), .B(B), .Y(n7));
endmodule

module operator_A_5 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_6 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n5), .Y(P));
sg13g2_o21ai_1 U2 (.A1(A), .A2(B), .B1(n3), .Y(n5));
sg13g2_inv_2 U3 (.A(n4), .Y(G));
sg13g2_nand2_2 U4 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U5 (.A(A), .B(B), .Y(n3));
endmodule

module operator_A_7 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_8 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_9 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_nand2_2 U3 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(G));
endmodule

module operator_A_10 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(B), .Y(n3));
sg13g2_xnor2_1 U2 (.A(A), .B(n3), .Y(P));
sg13g2_inv_2 U3 (.A(n4), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n4));
endmodule

module operator_A_11 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n3));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_xnor2_1 U4 (.A(A), .B(B), .Y(n4));
endmodule

module operator_A_12 (A, B, G, P);
input A, B;
output G, P;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n2));
sg13g2_inv_2 U2 (.A(A), .Y(n1));
sg13g2_xnor2_1 U3 (.A(B), .B(n1), .Y(P));
sg13g2_inv_2 U4 (.A(n2), .Y(G));
endmodule

module operator_A_13 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n5), .Y(G));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n5));
sg13g2_inv_2 U3 (.A(A), .Y(n3));
sg13g2_inv_2 U4 (.A(B), .Y(n4));
sg13g2_nand2_2 U5 (.A(n3), .B(n4), .Y(n6));
sg13g2_nand2_2 U6 (.A(n5), .B(n6), .Y(n7));
sg13g2_inv_2 U7 (.A(n7), .Y(P));
endmodule

module operator_A_14 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_xnor2_1 U4 (.A(A), .B(B), .Y(n4));
endmodule

module operator_A_15 (A, B, G, P);
input A, B;
output G, P;

sg13g2_nand2_2 U1 (.A(n3), .B(n4), .Y(n5));
sg13g2_nand2_2 U2 (.A(n6), .B(n5), .Y(n7));
sg13g2_inv_2 U3 (.A(A), .Y(n3));
sg13g2_inv_2 U4 (.A(B), .Y(n4));
sg13g2_inv_2 U5 (.A(n6), .Y(G));
sg13g2_inv_2 U6 (.A(n7), .Y(P));
sg13g2_nand2_2 U7 (.A(A), .B(B), .Y(n6));
endmodule

module operator_A_16 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(n1), .B(B), .Y(P));
sg13g2_inv_2 U2 (.A(A), .Y(n1));
sg13g2_nand2_2 U3 (.A(B), .B(A), .Y(n2));
sg13g2_inv_2 U4 (.A(n2), .Y(G));
endmodule

module operator_A_17 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(B), .B(A), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(P));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_18 (A, B, G, P);
input A, B;
output G, P;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n5));
sg13g2_nand2_2 U2 (.A(n3), .B(n4), .Y(n6));
sg13g2_nand2_2 U3 (.A(n5), .B(n6), .Y(n8));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n7));
sg13g2_inv_2 U5 (.A(B), .Y(n3));
sg13g2_inv_2 U6 (.A(A), .Y(n4));
sg13g2_inv_2 U7 (.A(n7), .Y(G));
sg13g2_inv_2 U8 (.A(n8), .Y(P));
endmodule

module operator_A_19 (A, B, G, P);
input A, B;
output G, P;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(G));
sg13g2_xnor2_1 U3 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U4 (.A(n4), .Y(P));
endmodule

module operator_A_20 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(P));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_21 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n3));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_xnor2_1 U4 (.A(B), .B(A), .Y(n4));
endmodule

module operator_A_22 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_23 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_24 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(B), .B(A), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_25 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_26 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_27 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n3), .Y(G));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(P));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_28 (A, B, G, P);
input A, B;
output G, P;

sg13g2_xnor2_1 U1 (.A(A), .B(n3), .Y(P));
sg13g2_inv_2 U2 (.A(B), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n4));
endmodule

module operator_A_29 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_30 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_31 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_A_32 (A, B, G, P);
input A, B;
output G, P;

sg13g2_inv_2 U1 (.A(n4), .Y(P));
sg13g2_xnor2_1 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(G));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n3));
endmodule

module operator_B_1 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_2 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U3 (.A(n1), .Y(Po));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_3 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_4 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n1));
sg13g2_nand2_2 U2 (.A(n2), .B(n3), .Y(Go));
sg13g2_inv_2 U3 (.A(G), .Y(n2));
sg13g2_nand2_2 U4 (.A(P), .B(G1), .Y(n3));
sg13g2_inv_2 U5 (.A(n1), .Y(Po));
endmodule

module operator_B_5 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n1), .Y(Po));
sg13g2_inv_2 U2 (.A(G), .Y(n2));
sg13g2_nand2_2 U3 (.A(P), .B(P1), .Y(n1));
sg13g2_nand2_2 U4 (.A(n2), .B(n3), .Y(Go));
sg13g2_nand2_2 U5 (.A(G1), .B(P), .Y(n3));
endmodule

module operator_B_6 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U3 (.A(n1), .Y(Po));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_7 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n1));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n1), .Y(Po));
endmodule

module operator_B_8 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n5));
sg13g2_inv_2 U2 (.A(n5), .Y(Po));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n4));
sg13g2_inv_2 U4 (.A(n4), .Y(Go));
endmodule

module operator_B_9 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_10 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n4));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n5));
sg13g2_inv_2 U4 (.A(n5), .Y(Po));
endmodule

module operator_B_11 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_12 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_13 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U4 (.A(n1), .Y(Po));
endmodule

module operator_B_14 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n1), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n1));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_15 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_nand2_2 U3 (.A(P), .B(P1), .Y(n1));
sg13g2_inv_2 U4 (.A(n1), .Y(Po));
endmodule

module operator_B_16 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_17 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_18 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_19 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_20 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_21 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_22 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n4));
sg13g2_inv_2 U3 (.A(n5), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n5));
endmodule

module operator_B_23 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P), .B(P1), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(P), .A2(G1), .B1(G), .Y(n3));
endmodule

module operator_B_24 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_25 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_26 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n1), .Y(Po));
endmodule

module operator_B_27 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(Po));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_28 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_nand2_2 U3 (.A(P), .B(P1), .Y(n1));
sg13g2_inv_2 U4 (.A(n1), .Y(Po));
endmodule

module operator_B_29 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_inv_2 U4 (.A(n4), .Y(Po));
endmodule

module operator_B_30 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U3 (.A1(P), .A2(G1), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_31 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_nand2_2 U1 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_32 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_33 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_34 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_35 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_36 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_37 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_38 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_39 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_nand2_2 U2 (.A(P), .B(P1), .Y(n4));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_a21oi_2 U4 (.A1(P), .A2(G1), .B1(G), .Y(n3));
endmodule

module operator_B_40 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n1), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n1));
sg13g2_a21oi_2 U3 (.A1(P), .A2(G1), .B1(G), .Y(n3));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_41 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n5), .Y(Po));
sg13g2_nand2_2 U2 (.A(P), .B(P1), .Y(n5));
sg13g2_inv_2 U3 (.A(n4), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(P), .A2(G1), .B1(G), .Y(n4));
endmodule

module operator_B_42 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n1), .Y(Po));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_nand2_2 U4 (.A(P), .B(P1), .Y(n1));
endmodule

module operator_B_43 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_44 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n3));
sg13g2_inv_2 U2 (.A(n4), .Y(Po));
sg13g2_nand2_2 U3 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U4 (.A(n3), .Y(Go));
endmodule

module operator_B_45 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_inv_2 U2 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U3 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_46 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_47 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n3));
sg13g2_inv_2 U3 (.A(n4), .Y(Po));
sg13g2_nand2_2 U4 (.A(P1), .B(P), .Y(n4));
endmodule

module operator_B_48 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_B_49 (G, G1, Go, P, P1, Po);
input G, G1, P, P1;
output Go, Po;

sg13g2_inv_2 U1 (.A(n4), .Y(Po));
sg13g2_nand2_2 U2 (.A(P1), .B(P), .Y(n4));
sg13g2_inv_2 U3 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U4 (.A1(G1), .A2(P), .B1(G), .Y(n3));
endmodule

module operator_C_1 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_2 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_3 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_4 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_5 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_6 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_7 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(G1), .A2(P), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_8 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_9 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_10 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n3), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n3));
endmodule

module operator_C_11 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_12 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_13 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_14 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_15 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_16 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_17 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_18 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_19 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_20 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_21 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_22 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_23 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_24 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_25 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_26 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_27 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_nor2_2 U1 (.A(n4), .B(G), .Y(n5));
sg13g2_inv_2 U2 (.A(n5), .Y(Go));
sg13g2_nor2_2 U3 (.A(n2), .B(n3), .Y(n4));
sg13g2_inv_2 U4 (.A(P), .Y(n2));
sg13g2_inv_2 U5 (.A(G1), .Y(n3));
endmodule

module operator_C_28 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_29 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(G1), .A2(P), .B1(G), .Y(n2));
endmodule

module operator_C_30 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module operator_C_31 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_a21oi_2 U1 (.A1(P), .A2(G1), .B1(G), .Y(n2));
sg13g2_inv_2 U2 (.A(n2), .Y(Go));
endmodule

module operator_C_32 (G, G1, Go, P);
input G, G1, P;
output Go;

sg13g2_inv_2 U1 (.A(n2), .Y(Go));
sg13g2_a21oi_2 U2 (.A1(P), .A2(G1), .B1(G), .Y(n2));
endmodule

module booth_array (\double[0], \double[1], \double[2], \double[3], \double[4], \double[5], \double[6], \double[7], \multiplier[0], \multiplier[1], \multiplier[2], \multiplier[3], \multiplier[4], \multiplier[5], \multiplier[6], \multiplier[7], \multiplier[8], \multiplier[9], \multiplier[10], \multiplier[11], \multiplier[12], \multiplier[13], \multiplier[14], \multiplier[15], \negation[0], \negation[1], \negation[2], \negation[3], \negation[4], \negation[5], \negation[6], \negation[7], \zero[0], \zero[1], \zero[2], \zero[3], \zero[4], \zero[5], \zero[6], \zero[7]);
input \multiplier[0], \multiplier[1], \multiplier[2], \multiplier[3], \multiplier[4], \multiplier[5], \multiplier[6], \multiplier[7], \multiplier[8], \multiplier[9], \multiplier[10], \multiplier[11], \multiplier[12], \multiplier[13], \multiplier[14], \multiplier[15];
output \double[0], \double[1], \double[2], \double[3], \double[4], \double[5], \double[6], \double[7], \negation[0], \negation[1], \negation[2], \negation[3], \negation[4], \negation[5], \negation[6], \negation[7], \zero[0], \zero[1], \zero[2], \zero[3], \zero[4], \zero[5], \zero[6], \zero[7];

sg13g2_inv_2 U2 (.A(n7), .Y(n1));
sg13g2_inv_2 U3 (.A(n1), .Y(\negation[7]));
sg13g2_inv_2 U4 (.A(n9), .Y(n5));
sg13g2_inv_2 U5 (.A(n5), .Y(\negation[2]));
sg13g2_inv_2 U6 (.A(n8), .Y(n3));
sg13g2_inv_2 U7 (.A(n3), .Y(\negation[3]));
sg13g2_tielo U8 (.L_LO(\*Logic0*));
booth_radix4_0 booth_radix4_0(.\codes[0](\*Logic0*), .\codes[1](\multiplier[0]), .\codes[2](\multiplier[1]), .double(\double[0]), .negation(\negation[0]), .zero(\zero[0]));
booth_radix4_1 booth_radix4_7(.\codes[0](\multiplier[13]), .\codes[1](\multiplier[14]), .\codes[2](\multiplier[15]), .double(\double[7]), .negation(n7), .zero(\zero[7]));
booth_radix4_2 booth_radix4_6(.\codes[0](\multiplier[11]), .\codes[1](\multiplier[12]), .\codes[2](\multiplier[13]), .double(\double[6]), .negation(\negation[6]), .zero(\zero[6]));
booth_radix4_3 booth_radix4_5(.\codes[0](\multiplier[9]), .\codes[1](\multiplier[10]), .\codes[2](\multiplier[11]), .double(\double[5]), .negation(\negation[5]), .zero(\zero[5]));
booth_radix4_4 booth_radix4_4(.\codes[0](\multiplier[7]), .\codes[1](\multiplier[8]), .\codes[2](\multiplier[9]), .double(\double[4]), .negation(\negation[4]), .zero(\zero[4]));
booth_radix4_5 booth_radix4_3(.\codes[0](\multiplier[5]), .\codes[1](\multiplier[6]), .\codes[2](\multiplier[7]), .double(\double[3]), .negation(n8), .zero(\zero[3]));
booth_radix4_6 booth_radix4_2(.\codes[0](\multiplier[3]), .\codes[1](\multiplier[4]), .\codes[2](\multiplier[5]), .double(\double[2]), .negation(n9), .zero(\zero[2]));
booth_radix4_7 booth_radix4_1(.\codes[0](\multiplier[1]), .\codes[1](\multiplier[2]), .\codes[2](\multiplier[3]), .double(\double[1]), .negation(\negation[1]), .zero(\zero[1]));
endmodule

module booth_radix4_0 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_nand3_1 U1 (.A(n1), .B(n4), .C(n5), .Y(n3));
sg13g2_nand3_1 U2 (.A(n1), .B(\codes[0]), .C(\codes[1]), .Y(n6));
sg13g2_nand2_2 U3 (.A(\codes[1]), .B(\codes[0]), .Y(n2));
sg13g2_nand3_1 U4 (.A(\codes[2]), .B(n4), .C(n5), .Y(n7));
sg13g2_nand2_2 U5 (.A(n6), .B(n7), .Y(double));
sg13g2_o21ai_1 U6 (.A1(n2), .A2(n1), .B1(n3), .Y(zero));
sg13g2_inv_2 U7 (.A(\codes[1]), .Y(n4));
sg13g2_inv_2 U8 (.A(\codes[0]), .Y(n5));
sg13g2_inv_2 U9 (.A(\codes[2]), .Y(n1));
sg13g2_a21oi_2 U10 (.A1(\codes[1]), .A2(\codes[0]), .B1(n1), .Y(negation));
endmodule

module booth_radix4_1 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_a21oi_2 U1 (.A1(\codes[1]), .A2(\codes[0]), .B1(n14), .Y(negation));
sg13g2_nand3_1 U2 (.A(n11), .B(n14), .C(n10), .Y(n12));
sg13g2_nand2_2 U3 (.A(\codes[1]), .B(\codes[0]), .Y(n13));
sg13g2_o21ai_1 U4 (.A1(n14), .A2(n13), .B1(n12), .Y(zero));
sg13g2_inv_2 U5 (.A(\codes[0]), .Y(n10));
sg13g2_nand3_1 U6 (.A(n10), .B(n11), .C(\codes[2]), .Y(n8));
sg13g2_inv_2 U7 (.A(\codes[1]), .Y(n11));
sg13g2_nand2_2 U8 (.A(n9), .B(n8), .Y(double));
sg13g2_nand3_1 U9 (.A(\codes[0]), .B(n14), .C(\codes[1]), .Y(n9));
sg13g2_inv_2 U10 (.A(\codes[2]), .Y(n14));
endmodule

module booth_radix4_2 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_nand3_1 U1 (.A(n10), .B(n11), .C(\codes[2]), .Y(n8));
sg13g2_nand3_1 U2 (.A(\codes[0]), .B(n14), .C(\codes[1]), .Y(n9));
sg13g2_nand2_2 U3 (.A(\codes[1]), .B(\codes[0]), .Y(n13));
sg13g2_inv_2 U4 (.A(\codes[0]), .Y(n10));
sg13g2_o21ai_1 U5 (.A1(n14), .A2(n13), .B1(n12), .Y(zero));
sg13g2_nand2_2 U6 (.A(n8), .B(n9), .Y(double));
sg13g2_inv_2 U7 (.A(\codes[1]), .Y(n11));
sg13g2_a21oi_2 U8 (.A1(\codes[1]), .A2(\codes[0]), .B1(n14), .Y(negation));
sg13g2_nand3_1 U9 (.A(n11), .B(n14), .C(n10), .Y(n12));
sg13g2_inv_2 U10 (.A(\codes[2]), .Y(n14));
endmodule

module booth_radix4_3 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_inv_2 U1 (.A(\codes[1]), .Y(n11));
sg13g2_nand3_1 U2 (.A(\codes[0]), .B(n14), .C(\codes[1]), .Y(n9));
sg13g2_nand3_1 U3 (.A(n10), .B(n11), .C(\codes[2]), .Y(n8));
sg13g2_a21oi_2 U4 (.A1(\codes[0]), .A2(\codes[1]), .B1(n14), .Y(negation));
sg13g2_nand2_2 U5 (.A(\codes[1]), .B(\codes[0]), .Y(n13));
sg13g2_inv_2 U6 (.A(\codes[0]), .Y(n10));
sg13g2_inv_2 U7 (.A(\codes[2]), .Y(n14));
sg13g2_nand2_2 U8 (.A(n9), .B(n8), .Y(double));
sg13g2_o21ai_1 U9 (.A1(n14), .A2(n13), .B1(n12), .Y(zero));
sg13g2_nand3_1 U10 (.A(n11), .B(n14), .C(n10), .Y(n12));
endmodule

module booth_radix4_4 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_inv_2 U1 (.A(n16), .Y(n9));
sg13g2_nand3_1 U2 (.A(n9), .B(n13), .C(n12), .Y(n10));
sg13g2_nand2_2 U3 (.A(\codes[0]), .B(\codes[1]), .Y(n15));
sg13g2_inv_2 U4 (.A(\codes[2]), .Y(n8));
sg13g2_nand3_1 U5 (.A(n16), .B(\codes[0]), .C(\codes[1]), .Y(n11));
sg13g2_o21ai_1 U6 (.A1(n8), .A2(n15), .B1(n14), .Y(zero));
sg13g2_nand3_1 U7 (.A(n12), .B(n16), .C(n13), .Y(n14));
sg13g2_inv_2 U8 (.A(\codes[1]), .Y(n13));
sg13g2_inv_2 U9 (.A(\codes[0]), .Y(n12));
sg13g2_nand2_2 U10 (.A(n11), .B(n10), .Y(double));
sg13g2_inv_2 U11 (.A(\codes[2]), .Y(n16));
sg13g2_a21oi_2 U12 (.A1(\codes[0]), .A2(\codes[1]), .B1(n16), .Y(negation));
endmodule

module booth_radix4_5 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_nand2_2 U1 (.A(n2), .B(n9), .Y(n4));
sg13g2_inv_2 U2 (.A(\codes[1]), .Y(n8));
sg13g2_nor2_2 U3 (.A(n8), .B(n14), .Y(n2));
sg13g2_nand3_1 U4 (.A(n14), .B(n12), .C(n8), .Y(n13));
sg13g2_nand3_1 U5 (.A(\codes[2]), .B(n12), .C(n8), .Y(n10));
sg13g2_inv_2 U6 (.A(\codes[0]), .Y(n12));
sg13g2_nand3_1 U7 (.A(n14), .B(n9), .C(\codes[1]), .Y(n11));
sg13g2_nand2_2 U8 (.A(n4), .B(n13), .Y(zero));
sg13g2_nand2_2 U9 (.A(n10), .B(n11), .Y(double));
sg13g2_inv_2 U10 (.A(\codes[2]), .Y(n14));
sg13g2_buf_2 U11 (.A(\codes[0]), .X(n9));
sg13g2_a21oi_2 U12 (.A1(\codes[0]), .A2(\codes[1]), .B1(n14), .Y(negation));
endmodule

module booth_radix4_6 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_buf_2 U1 (.A(\codes[2]), .X(n8));
sg13g2_nand2_2 U2 (.A(n8), .B(n9), .Y(n10));
sg13g2_nand2_2 U3 (.A(n10), .B(n15), .Y(zero));
sg13g2_inv_2 U4 (.A(n16), .Y(n9));
sg13g2_nand2_2 U5 (.A(\codes[0]), .B(\codes[1]), .Y(n16));
sg13g2_nand3_1 U6 (.A(\codes[0]), .B(n17), .C(\codes[1]), .Y(n12));
sg13g2_inv_2 U7 (.A(\codes[1]), .Y(n14));
sg13g2_nand3_1 U8 (.A(n8), .B(n13), .C(n14), .Y(n11));
sg13g2_inv_2 U9 (.A(\codes[0]), .Y(n13));
sg13g2_nand3_1 U10 (.A(n13), .B(n17), .C(n14), .Y(n15));
sg13g2_nand2_2 U11 (.A(n11), .B(n12), .Y(double));
sg13g2_a21oi_2 U12 (.A1(\codes[0]), .A2(\codes[1]), .B1(n17), .Y(negation));
sg13g2_inv_2 U13 (.A(\codes[2]), .Y(n17));
endmodule

module booth_radix4_7 (\codes[0], \codes[1], \codes[2], double, negation, zero);
input \codes[0], \codes[1], \codes[2];
output double, negation, zero;

sg13g2_inv_2 U1 (.A(\codes[2]), .Y(n14));
sg13g2_nand3_1 U2 (.A(\codes[0]), .B(n14), .C(\codes[1]), .Y(n9));
sg13g2_nand2_2 U3 (.A(\codes[0]), .B(\codes[1]), .Y(n13));
sg13g2_nand3_1 U4 (.A(n14), .B(n11), .C(n10), .Y(n12));
sg13g2_o21ai_1 U5 (.A1(n14), .A2(n13), .B1(n12), .Y(zero));
sg13g2_nand3_1 U6 (.A(\codes[2]), .B(n10), .C(n11), .Y(n8));
sg13g2_inv_2 U7 (.A(\codes[0]), .Y(n10));
sg13g2_inv_2 U8 (.A(\codes[1]), .Y(n11));
sg13g2_a21oi_2 U9 (.A1(\codes[0]), .A2(\codes[1]), .B1(n14), .Y(negation));
sg13g2_nand2_2 U10 (.A(n8), .B(n9), .Y(double));
endmodule

module compressor42_0 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n1), .B(n2), .Y(cout));
sg13g2_xnor2_1 U2 (.A(n4), .B(n3), .Y(n9));
sg13g2_inv_2 U3 (.A(n6), .Y(n5));
sg13g2_o21ai_1 U4 (.A1(D), .A2(C), .B1(n1), .Y(n4));
sg13g2_o21ai_1 U5 (.A1(A), .A2(B), .B1(n2), .Y(n3));
sg13g2_nand2_2 U6 (.A(n8), .B(cin), .Y(n7));
sg13g2_xnor2_1 U7 (.A(n9), .B(cin), .Y(S));
sg13g2_buf_2 U8 (.A(n4), .X(n10));
sg13g2_inv_2 U9 (.A(n9), .Y(n8));
sg13g2_o21ai_1 U10 (.A1(n10), .A2(n11), .B1(n5), .Y(carry));
sg13g2_o21ai_1 U11 (.A1(A), .A2(B), .B1(n2), .Y(n11));
sg13g2_nand2_2 U12 (.A(B), .B(A), .Y(n2));
sg13g2_o21ai_1 U13 (.A1(n1), .A2(n2), .B1(n7), .Y(n6));
sg13g2_nand2_2 U14 (.A(C), .B(D), .Y(n1));
endmodule

module compressor42_1 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n30), .B(n31), .Y(cout));
sg13g2_inv_2 U2 (.A(C), .Y(n15));
sg13g2_nand2_2 U3 (.A(C), .B(D), .Y(n31));
sg13g2_nand2_2 U4 (.A(n19), .B(n30), .Y(n10));
sg13g2_nand2_2 U5 (.A(A), .B(B), .Y(n30));
sg13g2_nand2_2 U6 (.A(n11), .B(n12), .Y(n13));
sg13g2_xnor2_1 U7 (.A(n23), .B(cin), .Y(S));
sg13g2_nand2_2 U8 (.A(n27), .B(n13), .Y(carry));
sg13g2_inv_2 U9 (.A(n10), .Y(n11));
sg13g2_inv_2 U10 (.A(n28), .Y(n12));
sg13g2_inv_2 U11 (.A(n26), .Y(n27));
sg13g2_nand2_2 U12 (.A(n15), .B(n14), .Y(n16));
sg13g2_nand2_2 U13 (.A(n16), .B(n31), .Y(n28));
sg13g2_inv_2 U14 (.A(D), .Y(n14));
sg13g2_nand2_2 U15 (.A(n25), .B(n22), .Y(n26));
sg13g2_nand2_2 U16 (.A(n24), .B(cin), .Y(n25));
sg13g2_xnor2_1 U17 (.A(n29), .B(n28), .Y(n23));
sg13g2_nand2_2 U18 (.A(n18), .B(n17), .Y(n19));
sg13g2_inv_2 U19 (.A(A), .Y(n18));
sg13g2_nand2_2 U20 (.A(n19), .B(n30), .Y(n29));
sg13g2_inv_2 U21 (.A(B), .Y(n17));
sg13g2_inv_2 U22 (.A(n23), .Y(n24));
sg13g2_nand2_2 U23 (.A(n20), .B(n21), .Y(n22));
sg13g2_inv_2 U24 (.A(n31), .Y(n20));
sg13g2_inv_2 U25 (.A(n30), .Y(n21));
endmodule

module compressor42_2 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n5), .B(n21), .Y(cout));
sg13g2_buf_2 U2 (.A(n20), .X(n5));
sg13g2_nand2_2 U3 (.A(n13), .B(n21), .Y(n6));
sg13g2_nor2_2 U4 (.A(n21), .B(n5), .Y(n9));
sg13g2_inv_2 U5 (.A(n9), .Y(n14));
sg13g2_inv_2 U6 (.A(n15), .Y(n16));
sg13g2_xnor2_1 U7 (.A(n15), .B(cin), .Y(S));
sg13g2_nand3_1 U8 (.A(n1), .B(n14), .C(n17), .Y(carry));
sg13g2_o21ai_1 U9 (.A1(B), .A2(A), .B1(n5), .Y(n10));
sg13g2_inv_2 U10 (.A(D), .Y(n11));
sg13g2_nand2_2 U11 (.A(n11), .B(n12), .Y(n13));
sg13g2_nand2_2 U12 (.A(n13), .B(n21), .Y(n18));
sg13g2_inv_2 U13 (.A(C), .Y(n12));
sg13g2_nand2_2 U14 (.A(n16), .B(cin), .Y(n17));
sg13g2_nand2_2 U15 (.A(D), .B(C), .Y(n21));
sg13g2_xnor2_1 U16 (.A(n18), .B(n19), .Y(n15));
sg13g2_o21ai_1 U17 (.A1(B), .A2(A), .B1(n20), .Y(n19));
sg13g2_nand2_2 U18 (.A(A), .B(B), .Y(n20));
sg13g2_or2_1 U19 (.A(n6), .B(n10), .X(n1));
endmodule

module compressor42_3 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n5), .B(n6), .Y(cout));
sg13g2_inv_2 U2 (.A(n14), .Y(n5));
sg13g2_buf_2 U3 (.A(n22), .X(n6));
sg13g2_nand2_2 U4 (.A(n10), .B(n11), .Y(n12));
sg13g2_nand3_1 U5 (.A(n15), .B(n1), .C(n18), .Y(carry));
sg13g2_inv_2 U6 (.A(n6), .Y(n13));
sg13g2_xnor2_1 U7 (.A(n16), .B(cin), .Y(S));
sg13g2_inv_2 U8 (.A(D), .Y(n10));
sg13g2_nand2_2 U9 (.A(D), .B(C), .Y(n22));
sg13g2_inv_2 U10 (.A(C), .Y(n11));
sg13g2_nand2_2 U11 (.A(n17), .B(cin), .Y(n18));
sg13g2_nand2_2 U12 (.A(n12), .B(n22), .Y(n19));
sg13g2_xnor2_1 U13 (.A(n19), .B(n20), .Y(n16));
sg13g2_nand2_2 U14 (.A(n13), .B(n14), .Y(n15));
sg13g2_inv_2 U15 (.A(n21), .Y(n14));
sg13g2_inv_2 U16 (.A(n16), .Y(n17));
sg13g2_o21ai_1 U17 (.A1(B), .A2(A), .B1(n21), .Y(n20));
sg13g2_nand2_2 U18 (.A(A), .B(B), .Y(n21));
sg13g2_or2_1 U19 (.A(n19), .B(n20), .X(n1));
endmodule

module compressor42_4 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n5), .B(n21), .Y(cout));
sg13g2_buf_2 U2 (.A(n20), .X(n5));
sg13g2_o21ai_1 U3 (.A1(C), .A2(D), .B1(n21), .Y(n18));
sg13g2_xnor2_1 U4 (.A(n19), .B(n18), .Y(n15));
sg13g2_nand2_2 U5 (.A(n16), .B(cin), .Y(n17));
sg13g2_inv_2 U6 (.A(n15), .Y(n16));
sg13g2_xnor2_1 U7 (.A(n15), .B(cin), .Y(S));
sg13g2_nand3_1 U8 (.A(n14), .B(n1), .C(n17), .Y(carry));
sg13g2_inv_2 U9 (.A(A), .Y(n10));
sg13g2_nand2_2 U10 (.A(D), .B(C), .Y(n21));
sg13g2_nand2_2 U11 (.A(n10), .B(n6), .Y(n11));
sg13g2_nand2_2 U12 (.A(n11), .B(n20), .Y(n19));
sg13g2_inv_2 U13 (.A(B), .Y(n6));
sg13g2_nand2_2 U14 (.A(n12), .B(n13), .Y(n14));
sg13g2_inv_2 U15 (.A(n21), .Y(n12));
sg13g2_inv_2 U16 (.A(n5), .Y(n13));
sg13g2_nand2_2 U17 (.A(A), .B(B), .Y(n20));
sg13g2_or2_1 U18 (.A(n19), .B(n18), .X(n1));
endmodule

module compressor42_5 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n16), .B(n15), .Y(cout));
sg13g2_inv_2 U2 (.A(n10), .Y(n11));
sg13g2_nor2_2 U3 (.A(n16), .B(n15), .Y(n5));
sg13g2_inv_2 U4 (.A(n5), .Y(n6));
sg13g2_nand2_2 U5 (.A(n11), .B(cin), .Y(n12));
sg13g2_nand3_1 U6 (.A(n1), .B(n6), .C(n12), .Y(carry));
sg13g2_xnor2_1 U7 (.A(n10), .B(cin), .Y(S));
sg13g2_o21ai_1 U8 (.A1(C), .A2(D), .B1(n16), .Y(n13));
sg13g2_nand2_2 U9 (.A(D), .B(C), .Y(n16));
sg13g2_xnor2_1 U10 (.A(n13), .B(n14), .Y(n10));
sg13g2_o21ai_1 U11 (.A1(B), .A2(A), .B1(n15), .Y(n14));
sg13g2_nand2_2 U12 (.A(A), .B(B), .Y(n15));
sg13g2_or2_1 U13 (.A(n14), .B(n13), .X(n1));
endmodule

module compressor42_6 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n28), .B(n29), .Y(cout));
sg13g2_buf_2 U2 (.A(n28), .X(n10));
sg13g2_o21ai_1 U3 (.A1(D), .A2(C), .B1(n29), .Y(n26));
sg13g2_inv_2 U4 (.A(n24), .Y(n25));
sg13g2_nand2_2 U5 (.A(n20), .B(n10), .Y(n11));
sg13g2_nand2_2 U6 (.A(n19), .B(n18), .Y(n20));
sg13g2_inv_2 U7 (.A(A), .Y(n19));
sg13g2_nand2_2 U8 (.A(A), .B(B), .Y(n28));
sg13g2_nand2_2 U9 (.A(n25), .B(n17), .Y(carry));
sg13g2_xnor2_1 U10 (.A(n21), .B(cin), .Y(S));
sg13g2_nand2_2 U11 (.A(n12), .B(n13), .Y(n14));
sg13g2_nand2_2 U12 (.A(n23), .B(n14), .Y(n24));
sg13g2_inv_2 U13 (.A(n29), .Y(n12));
sg13g2_inv_2 U14 (.A(n10), .Y(n13));
sg13g2_nand2_2 U15 (.A(C), .B(D), .Y(n29));
sg13g2_xnor2_1 U16 (.A(n26), .B(n27), .Y(n21));
sg13g2_nand2_2 U17 (.A(n22), .B(cin), .Y(n23));
sg13g2_inv_2 U18 (.A(n21), .Y(n22));
sg13g2_nand2_2 U19 (.A(n15), .B(n16), .Y(n17));
sg13g2_inv_2 U20 (.A(n11), .Y(n15));
sg13g2_inv_2 U21 (.A(n26), .Y(n16));
sg13g2_nand2_2 U22 (.A(n20), .B(n28), .Y(n27));
sg13g2_inv_2 U23 (.A(B), .Y(n18));
endmodule

module compressor42_7 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n8), .B(n31), .Y(cout));
sg13g2_buf_2 U2 (.A(n30), .X(n8));
sg13g2_o21ai_1 U3 (.A1(A), .A2(B), .B1(n30), .Y(n29));
sg13g2_nand2_2 U4 (.A(n20), .B(n31), .Y(n10));
sg13g2_inv_2 U5 (.A(C), .Y(n19));
sg13g2_nand2_2 U6 (.A(n11), .B(cin), .Y(n25));
sg13g2_nand2_2 U7 (.A(n11), .B(n12), .Y(n14));
sg13g2_nand2_2 U8 (.A(n13), .B(n14), .Y(S));
sg13g2_inv_2 U9 (.A(n24), .Y(n11));
sg13g2_nand2_2 U10 (.A(n24), .B(cin), .Y(n13));
sg13g2_inv_2 U11 (.A(cin), .Y(n12));
sg13g2_xnor2_1 U12 (.A(n29), .B(n28), .Y(n24));
sg13g2_nand2_2 U13 (.A(n15), .B(n16), .Y(n17));
sg13g2_nand2_2 U14 (.A(n27), .B(n17), .Y(carry));
sg13g2_inv_2 U15 (.A(n29), .Y(n15));
sg13g2_inv_2 U16 (.A(n10), .Y(n16));
sg13g2_inv_2 U17 (.A(n26), .Y(n27));
sg13g2_nand2_2 U18 (.A(n18), .B(n19), .Y(n20));
sg13g2_nand2_2 U19 (.A(n20), .B(n31), .Y(n28));
sg13g2_inv_2 U20 (.A(D), .Y(n18));
sg13g2_nand2_2 U21 (.A(D), .B(C), .Y(n31));
sg13g2_nand2_2 U22 (.A(A), .B(B), .Y(n30));
sg13g2_nand2_2 U23 (.A(n25), .B(n23), .Y(n26));
sg13g2_nand2_2 U24 (.A(n21), .B(n22), .Y(n23));
sg13g2_inv_2 U25 (.A(n31), .Y(n21));
sg13g2_inv_2 U26 (.A(n8), .Y(n22));
endmodule

module compressor42_8 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n14), .B(n24), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n15));
sg13g2_xnor2_1 U3 (.A(n23), .B(n22), .Y(n20));
sg13g2_nand3_1 U4 (.A(n8), .B(n1), .C(n21), .Y(carry));
sg13g2_o21ai_1 U5 (.A1(A), .A2(B), .B1(n15), .Y(n2));
sg13g2_inv_2 U6 (.A(n2), .Y(n6));
sg13g2_nand2_2 U7 (.A(n19), .B(n24), .Y(n5));
sg13g2_xnor2_1 U8 (.A(cin), .B(n20), .Y(S));
sg13g2_nand2_2 U9 (.A(n6), .B(n13), .Y(n8));
sg13g2_inv_2 U10 (.A(n20), .Y(n16));
sg13g2_nand2_2 U11 (.A(n10), .B(n11), .Y(n12));
sg13g2_nand2_2 U12 (.A(n12), .B(n15), .Y(n23));
sg13g2_inv_2 U13 (.A(A), .Y(n10));
sg13g2_inv_2 U14 (.A(B), .Y(n11));
sg13g2_inv_2 U15 (.A(n5), .Y(n13));
sg13g2_nand2_2 U16 (.A(A), .B(B), .Y(n14));
sg13g2_nand2_2 U17 (.A(n17), .B(n18), .Y(n19));
sg13g2_nand2_2 U18 (.A(D), .B(C), .Y(n24));
sg13g2_inv_2 U19 (.A(C), .Y(n18));
sg13g2_nand2_2 U20 (.A(n16), .B(cin), .Y(n21));
sg13g2_nand2_2 U21 (.A(n19), .B(n24), .Y(n22));
sg13g2_inv_2 U22 (.A(D), .Y(n17));
sg13g2_or2_1 U23 (.A(n24), .B(n14), .X(n1));
endmodule

module compressor42_9 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n17), .B(n16), .Y(cout));
sg13g2_nand3_1 U2 (.A(n13), .B(n1), .C(n10), .Y(carry));
sg13g2_o21ai_1 U3 (.A1(B), .A2(A), .B1(n16), .Y(n15));
sg13g2_nand2_2 U4 (.A(n12), .B(cin), .Y(n13));
sg13g2_xnor2_1 U5 (.A(n15), .B(n14), .Y(n11));
sg13g2_inv_2 U6 (.A(n11), .Y(n12));
sg13g2_xnor2_1 U7 (.A(n11), .B(cin), .Y(S));
sg13g2_o21ai_1 U8 (.A1(D), .A2(C), .B1(n17), .Y(n14));
sg13g2_nand2_2 U9 (.A(D), .B(C), .Y(n17));
sg13g2_nand2_2 U10 (.A(n5), .B(n6), .Y(n10));
sg13g2_inv_2 U11 (.A(n17), .Y(n5));
sg13g2_inv_2 U12 (.A(n16), .Y(n6));
sg13g2_nand2_2 U13 (.A(B), .B(A), .Y(n16));
sg13g2_or2_1 U14 (.A(n15), .B(n14), .X(n1));
endmodule

module compressor42_10 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n23), .B(n22), .Y(cout));
sg13g2_nand3_1 U2 (.A(n19), .B(n10), .C(n16), .Y(carry));
sg13g2_nand2_2 U3 (.A(n13), .B(n23), .Y(n20));
sg13g2_nand2_2 U4 (.A(C), .B(D), .Y(n23));
sg13g2_nand2_2 U5 (.A(n5), .B(n6), .Y(n10));
sg13g2_inv_2 U6 (.A(n17), .Y(n18));
sg13g2_xnor2_1 U7 (.A(n17), .B(cin), .Y(S));
sg13g2_xnor2_1 U8 (.A(n21), .B(n20), .Y(n17));
sg13g2_inv_2 U9 (.A(n23), .Y(n5));
sg13g2_inv_2 U10 (.A(n22), .Y(n6));
sg13g2_o21ai_1 U11 (.A1(B), .A2(A), .B1(n22), .Y(n21));
sg13g2_nand2_2 U12 (.A(n18), .B(cin), .Y(n19));
sg13g2_nand2_2 U13 (.A(n11), .B(n12), .Y(n13));
sg13g2_inv_2 U14 (.A(D), .Y(n11));
sg13g2_inv_2 U15 (.A(C), .Y(n12));
sg13g2_nand2_2 U16 (.A(n14), .B(n15), .Y(n16));
sg13g2_inv_2 U17 (.A(n21), .Y(n14));
sg13g2_inv_2 U18 (.A(n20), .Y(n15));
sg13g2_nand2_2 U19 (.A(B), .B(A), .Y(n22));
endmodule

module compressor42_11 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n18), .B(n17), .Y(cout));
sg13g2_inv_2 U2 (.A(n13), .Y(n14));
sg13g2_o21ai_1 U3 (.A1(n18), .A2(n17), .B1(n12), .Y(n13));
sg13g2_nand2_2 U4 (.A(n11), .B(cin), .Y(n12));
sg13g2_inv_2 U5 (.A(n10), .Y(n11));
sg13g2_o21ai_1 U6 (.A1(D), .A2(C), .B1(n18), .Y(n15));
sg13g2_xnor2_1 U7 (.A(n10), .B(cin), .Y(S));
sg13g2_xnor2_1 U8 (.A(n15), .B(n16), .Y(n10));
sg13g2_nand2_2 U9 (.A(A), .B(B), .Y(n17));
sg13g2_o21ai_1 U10 (.A1(A), .A2(B), .B1(n17), .Y(n16));
sg13g2_o21ai_1 U11 (.A1(n16), .A2(n15), .B1(n14), .Y(carry));
sg13g2_nand2_2 U12 (.A(C), .B(D), .Y(n18));
endmodule

module compressor42_12 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n23), .B(n22), .Y(cout));
sg13g2_nand3_1 U2 (.A(n16), .B(n1), .C(n19), .Y(carry));
sg13g2_nand2_2 U3 (.A(C), .B(D), .Y(n23));
sg13g2_xnor2_1 U4 (.A(n21), .B(n20), .Y(n17));
sg13g2_inv_2 U5 (.A(B), .Y(n5));
sg13g2_inv_2 U6 (.A(C), .Y(n12));
sg13g2_xnor2_1 U7 (.A(n17), .B(cin), .Y(S));
sg13g2_nand2_2 U8 (.A(n5), .B(n6), .Y(n10));
sg13g2_inv_2 U9 (.A(A), .Y(n6));
sg13g2_nand2_2 U10 (.A(B), .B(A), .Y(n22));
sg13g2_inv_2 U11 (.A(n17), .Y(n18));
sg13g2_nand2_2 U12 (.A(n13), .B(n23), .Y(n20));
sg13g2_inv_2 U13 (.A(D), .Y(n11));
sg13g2_nand2_2 U14 (.A(n10), .B(n22), .Y(n21));
sg13g2_nand2_2 U15 (.A(n11), .B(n12), .Y(n13));
sg13g2_nand2_2 U16 (.A(n14), .B(n15), .Y(n16));
sg13g2_inv_2 U17 (.A(n23), .Y(n14));
sg13g2_inv_2 U18 (.A(n22), .Y(n15));
sg13g2_nand2_2 U19 (.A(n18), .B(cin), .Y(n19));
sg13g2_or2_1 U20 (.A(n21), .B(n20), .X(n1));
endmodule

module compressor42_13 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n28), .B(n29), .Y(cout));
sg13g2_buf_2 U2 (.A(n27), .X(n5));
sg13g2_nand2_2 U3 (.A(n19), .B(n29), .Y(n6));
sg13g2_inv_2 U4 (.A(C), .Y(n18));
sg13g2_nand3_1 U5 (.A(n25), .B(n1), .C(n13), .Y(carry));
sg13g2_or2_1 U6 (.A(n5), .B(n6), .X(n1));
sg13g2_nand2_2 U7 (.A(n24), .B(cin), .Y(n25));
sg13g2_nand2_2 U8 (.A(n23), .B(cin), .Y(n21));
sg13g2_inv_2 U9 (.A(n23), .Y(n24));
sg13g2_nand2_2 U10 (.A(C), .B(D), .Y(n29));
sg13g2_nand2_2 U11 (.A(n11), .B(n12), .Y(n13));
sg13g2_inv_2 U12 (.A(n29), .Y(n11));
sg13g2_inv_2 U13 (.A(n28), .Y(n12));
sg13g2_nand2_2 U14 (.A(B), .B(A), .Y(n28));
sg13g2_nand2_2 U15 (.A(n14), .B(n15), .Y(n16));
sg13g2_nand2_2 U16 (.A(n28), .B(n16), .Y(n27));
sg13g2_inv_2 U17 (.A(A), .Y(n14));
sg13g2_inv_2 U18 (.A(B), .Y(n15));
sg13g2_nand2_2 U19 (.A(n17), .B(n18), .Y(n19));
sg13g2_nand2_2 U20 (.A(n19), .B(n29), .Y(n26));
sg13g2_inv_2 U21 (.A(D), .Y(n17));
sg13g2_xnor2_1 U22 (.A(n27), .B(n26), .Y(n23));
sg13g2_nand2_2 U23 (.A(n24), .B(n20), .Y(n22));
sg13g2_nand2_2 U24 (.A(n22), .B(n21), .Y(S));
sg13g2_inv_2 U25 (.A(cin), .Y(n20));
endmodule

module compressor42_14 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n29), .B(n28), .Y(cout));
sg13g2_nand2_2 U2 (.A(n18), .B(n19), .Y(n20));
sg13g2_inv_2 U3 (.A(B), .Y(n19));
sg13g2_inv_2 U4 (.A(n28), .Y(n5));
sg13g2_nand3_1 U5 (.A(n12), .B(n1), .C(n25), .Y(carry));
sg13g2_inv_2 U6 (.A(n27), .Y(n9));
sg13g2_nand2_2 U7 (.A(n9), .B(n17), .Y(n12));
sg13g2_inv_2 U8 (.A(n18), .Y(n8));
sg13g2_inv_2 U9 (.A(A), .Y(n18));
sg13g2_nand2_2 U10 (.A(n27), .B(n17), .Y(n10));
sg13g2_nand2_2 U11 (.A(n16), .B(n13), .Y(n15));
sg13g2_nand2b_1 U12 (.A_N(n29), .B(n5), .Y(n1));
sg13g2_inv_2 U13 (.A(n26), .Y(n17));
sg13g2_inv_2 U14 (.A(n16), .Y(n24));
sg13g2_inv_2 U15 (.A(C), .Y(n22));
sg13g2_nand2_2 U16 (.A(n9), .B(n26), .Y(n11));
sg13g2_nand2_2 U17 (.A(n10), .B(n11), .Y(n16));
sg13g2_nand2_2 U18 (.A(n24), .B(cin), .Y(n14));
sg13g2_nand2_2 U19 (.A(n14), .B(n15), .Y(S));
sg13g2_inv_2 U20 (.A(cin), .Y(n13));
sg13g2_nand2_2 U21 (.A(n21), .B(n22), .Y(n23));
sg13g2_nand2_2 U22 (.A(n16), .B(cin), .Y(n25));
sg13g2_nand2_2 U23 (.A(C), .B(D), .Y(n29));
sg13g2_nand2_2 U24 (.A(n20), .B(n28), .Y(n27));
sg13g2_nand2_2 U25 (.A(n23), .B(n29), .Y(n26));
sg13g2_inv_2 U26 (.A(D), .Y(n21));
sg13g2_nand2_2 U27 (.A(B), .B(n8), .Y(n28));
endmodule

module compressor42_15 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_inv_2 U1 (.A(D), .Y(n20));
sg13g2_nand2_2 U2 (.A(n24), .B(n6), .Y(n11));
sg13g2_nand2_2 U3 (.A(n22), .B(n29), .Y(n5));
sg13g2_nand3_1 U4 (.A(n25), .B(n19), .C(n14), .Y(carry));
sg13g2_nand2_2 U5 (.A(D), .B(C), .Y(n29));
sg13g2_inv_2 U6 (.A(C), .Y(n21));
sg13g2_nand2_2 U7 (.A(A), .B(B), .Y(n15));
sg13g2_nand2_2 U8 (.A(n23), .B(cin), .Y(n10));
sg13g2_nand2_2 U9 (.A(n10), .B(n11), .Y(S));
sg13g2_inv_2 U10 (.A(cin), .Y(n6));
sg13g2_o21ai_1 U11 (.A1(B), .A2(A), .B1(n15), .Y(n12));
sg13g2_nand2_2 U12 (.A(n21), .B(n20), .Y(n22));
sg13g2_nand2_2 U13 (.A(n29), .B(n15), .Y(cout));
sg13g2_inv_2 U14 (.A(n29), .Y(n16));
sg13g2_xnor2_1 U15 (.A(n27), .B(n26), .Y(n23));
sg13g2_nand2_2 U16 (.A(n13), .B(n17), .Y(n14));
sg13g2_inv_2 U17 (.A(n12), .Y(n13));
sg13g2_nand2_2 U18 (.A(n24), .B(cin), .Y(n25));
sg13g2_o21ai_1 U19 (.A1(B), .A2(A), .B1(n28), .Y(n27));
sg13g2_inv_2 U20 (.A(n5), .Y(n17));
sg13g2_inv_2 U21 (.A(n23), .Y(n24));
sg13g2_nand2_2 U22 (.A(n16), .B(n18), .Y(n19));
sg13g2_inv_2 U23 (.A(n15), .Y(n18));
sg13g2_nand2_2 U24 (.A(n22), .B(n29), .Y(n26));
sg13g2_nand2_2 U25 (.A(A), .B(B), .Y(n28));
endmodule

module compressor42_16 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n28), .B(n27), .Y(cout));
sg13g2_nand3_1 U2 (.A(n24), .B(n10), .C(n14), .Y(carry));
sg13g2_inv_2 U3 (.A(n25), .Y(n11));
sg13g2_nand2_2 U4 (.A(n23), .B(cin), .Y(n24));
sg13g2_inv_2 U5 (.A(C), .Y(n19));
sg13g2_nand2_2 U6 (.A(n5), .B(n6), .Y(n10));
sg13g2_inv_2 U7 (.A(n28), .Y(n5));
sg13g2_inv_2 U8 (.A(n27), .Y(n6));
sg13g2_inv_2 U9 (.A(D), .Y(n20));
sg13g2_inv_2 U10 (.A(n26), .Y(n15));
sg13g2_xnor2_1 U11 (.A(n22), .B(cin), .Y(S));
sg13g2_nand2_2 U12 (.A(B), .B(A), .Y(n27));
sg13g2_nand2_2 U13 (.A(n25), .B(n26), .Y(n12));
sg13g2_nand2_2 U14 (.A(n15), .B(n11), .Y(n13));
sg13g2_nand2_2 U15 (.A(n13), .B(n12), .Y(n22));
sg13g2_inv_2 U16 (.A(n22), .Y(n23));
sg13g2_nand2_2 U17 (.A(n21), .B(n28), .Y(n25));
sg13g2_nand2_2 U18 (.A(n15), .B(n11), .Y(n14));
sg13g2_nand2_2 U19 (.A(n16), .B(n17), .Y(n18));
sg13g2_nand2_2 U20 (.A(n18), .B(n27), .Y(n26));
sg13g2_inv_2 U21 (.A(B), .Y(n16));
sg13g2_inv_2 U22 (.A(A), .Y(n17));
sg13g2_nand2_2 U23 (.A(n19), .B(n20), .Y(n21));
sg13g2_nand2_2 U24 (.A(D), .B(C), .Y(n28));
endmodule

module compressor42_17 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n11), .B(n23), .Y(cout));
sg13g2_xnor2_1 U2 (.A(n21), .B(n22), .Y(n18));
sg13g2_xnor2_1 U3 (.A(n18), .B(cin), .Y(S));
sg13g2_nand3_1 U4 (.A(n17), .B(n1), .C(n20), .Y(carry));
sg13g2_nand2_2 U5 (.A(n13), .B(n12), .Y(n5));
sg13g2_nand2_2 U6 (.A(n5), .B(n23), .Y(n6));
sg13g2_nand2_2 U7 (.A(D), .B(C), .Y(n24));
sg13g2_o21ai_1 U8 (.A1(C), .A2(D), .B1(n24), .Y(n10));
sg13g2_nand2_2 U9 (.A(B), .B(A), .Y(n23));
sg13g2_nand2_2 U10 (.A(D), .B(C), .Y(n11));
sg13g2_nand2_2 U11 (.A(n19), .B(cin), .Y(n20));
sg13g2_inv_2 U12 (.A(n18), .Y(n19));
sg13g2_inv_2 U13 (.A(B), .Y(n12));
sg13g2_nand2_2 U14 (.A(n12), .B(n13), .Y(n14));
sg13g2_nand2_2 U15 (.A(n14), .B(n23), .Y(n22));
sg13g2_inv_2 U16 (.A(A), .Y(n13));
sg13g2_nand2_2 U17 (.A(n15), .B(n16), .Y(n17));
sg13g2_inv_2 U18 (.A(n23), .Y(n15));
sg13g2_inv_2 U19 (.A(n11), .Y(n16));
sg13g2_o21ai_1 U20 (.A1(C), .A2(D), .B1(n24), .Y(n21));
sg13g2_or2_1 U21 (.A(n6), .B(n10), .X(n1));
endmodule

module compressor42_18 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n5), .B(n23), .Y(cout));
sg13g2_inv_2 U2 (.A(n12), .Y(n5));
sg13g2_inv_2 U3 (.A(n24), .Y(n12));
sg13g2_inv_2 U4 (.A(C), .Y(n16));
sg13g2_nand2_2 U5 (.A(n17), .B(n24), .Y(n6));
sg13g2_nor2_2 U6 (.A(n22), .B(n6), .Y(n10));
sg13g2_inv_2 U7 (.A(n10), .Y(n11));
sg13g2_o21ai_1 U8 (.A1(A), .A2(B), .B1(n23), .Y(n22));
sg13g2_nand3_1 U9 (.A(n14), .B(n20), .C(n11), .Y(carry));
sg13g2_nand2_2 U10 (.A(n19), .B(cin), .Y(n20));
sg13g2_inv_2 U11 (.A(D), .Y(n15));
sg13g2_xnor2_1 U12 (.A(n22), .B(n21), .Y(n18));
sg13g2_nand2_2 U13 (.A(n15), .B(n16), .Y(n17));
sg13g2_xnor2_1 U14 (.A(n18), .B(cin), .Y(S));
sg13g2_inv_2 U15 (.A(n18), .Y(n19));
sg13g2_inv_2 U16 (.A(n23), .Y(n13));
sg13g2_nand2_2 U17 (.A(n12), .B(n13), .Y(n14));
sg13g2_nand2_2 U18 (.A(B), .B(A), .Y(n23));
sg13g2_nand2_2 U19 (.A(n17), .B(n24), .Y(n21));
sg13g2_nand2_2 U20 (.A(D), .B(C), .Y(n24));
endmodule

module compressor42_19 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n27), .B(n26), .Y(cout));
sg13g2_inv_2 U2 (.A(D), .Y(n15));
sg13g2_xnor2_1 U3 (.A(n10), .B(cin), .Y(S));
sg13g2_nand3_1 U4 (.A(n20), .B(n1), .C(n23), .Y(carry));
sg13g2_nand2_2 U5 (.A(n14), .B(n26), .Y(n5));
sg13g2_nand2_2 U6 (.A(n14), .B(n26), .Y(n6));
sg13g2_nand2_2 U7 (.A(n12), .B(n13), .Y(n14));
sg13g2_xnor2_1 U8 (.A(n5), .B(n24), .Y(n10));
sg13g2_xnor2_1 U9 (.A(n25), .B(n24), .Y(n21));
sg13g2_nand2_2 U10 (.A(n17), .B(n27), .Y(n11));
sg13g2_inv_2 U11 (.A(A), .Y(n13));
sg13g2_nand2_2 U12 (.A(n22), .B(cin), .Y(n23));
sg13g2_nand2_2 U13 (.A(n14), .B(n26), .Y(n25));
sg13g2_inv_2 U14 (.A(B), .Y(n12));
sg13g2_inv_2 U15 (.A(n21), .Y(n22));
sg13g2_nand2_2 U16 (.A(n15), .B(n16), .Y(n17));
sg13g2_nand2_2 U17 (.A(n17), .B(n27), .Y(n24));
sg13g2_inv_2 U18 (.A(C), .Y(n16));
sg13g2_nand2_2 U19 (.A(n18), .B(n19), .Y(n20));
sg13g2_inv_2 U20 (.A(n27), .Y(n18));
sg13g2_inv_2 U21 (.A(n26), .Y(n19));
sg13g2_nand2_2 U22 (.A(B), .B(A), .Y(n26));
sg13g2_nand2_2 U23 (.A(C), .B(D), .Y(n27));
sg13g2_or2_1 U24 (.A(n11), .B(n6), .X(n1));
endmodule

module compressor42_20 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(D), .B(C), .Y(n30));
sg13g2_buf_2 U2 (.A(n30), .X(n10));
sg13g2_inv_2 U3 (.A(D), .Y(n15));
sg13g2_inv_2 U4 (.A(B), .Y(n19));
sg13g2_inv_2 U5 (.A(A), .Y(n20));
sg13g2_xnor2_1 U6 (.A(n12), .B(cin), .Y(S));
sg13g2_inv_2 U7 (.A(n23), .Y(n11));
sg13g2_xnor2_1 U8 (.A(n27), .B(n28), .Y(n22));
sg13g2_buf_2 U9 (.A(n11), .X(n12));
sg13g2_nand2_2 U10 (.A(n29), .B(n10), .Y(cout));
sg13g2_inv_2 U11 (.A(n27), .Y(n13));
sg13g2_o21ai_1 U12 (.A1(n10), .A2(n29), .B1(n24), .Y(n25));
sg13g2_nand2_2 U13 (.A(B), .B(A), .Y(n29));
sg13g2_nand2_2 U14 (.A(n14), .B(n15), .Y(n16));
sg13g2_nand2_2 U15 (.A(n16), .B(n30), .Y(n27));
sg13g2_inv_2 U16 (.A(C), .Y(n14));
sg13g2_nand2_2 U17 (.A(n17), .B(n13), .Y(n18));
sg13g2_nand2_2 U18 (.A(n26), .B(n18), .Y(carry));
sg13g2_inv_2 U19 (.A(n28), .Y(n17));
sg13g2_inv_2 U20 (.A(n25), .Y(n26));
sg13g2_nand2_2 U21 (.A(n23), .B(cin), .Y(n24));
sg13g2_inv_2 U22 (.A(n22), .Y(n23));
sg13g2_nand2_2 U23 (.A(n19), .B(n20), .Y(n21));
sg13g2_nand2_2 U24 (.A(n21), .B(n29), .Y(n28));
endmodule

module compressor42_21 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n20), .B(n19), .Y(cout));
sg13g2_inv_2 U2 (.A(n13), .Y(n10));
sg13g2_o21ai_1 U3 (.A1(B), .A2(A), .B1(n19), .Y(n18));
sg13g2_xnor2_1 U4 (.A(n18), .B(n17), .Y(n12));
sg13g2_xnor2_1 U5 (.A(n10), .B(cin), .Y(S));
sg13g2_nand2_2 U6 (.A(D), .B(C), .Y(n20));
sg13g2_o21ai_1 U7 (.A1(D), .A2(C), .B1(n20), .Y(n17));
sg13g2_o21ai_1 U8 (.A1(n11), .A2(n17), .B1(n16), .Y(carry));
sg13g2_inv_2 U9 (.A(n12), .Y(n13));
sg13g2_buf_2 U10 (.A(n18), .X(n11));
sg13g2_nand2_2 U11 (.A(B), .B(A), .Y(n19));
sg13g2_inv_2 U12 (.A(n15), .Y(n16));
sg13g2_o21ai_1 U13 (.A1(n19), .A2(n20), .B1(n14), .Y(n15));
sg13g2_nand2_2 U14 (.A(n13), .B(cin), .Y(n14));
endmodule

module compressor42_22 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n19), .B(n20), .Y(cout));
sg13g2_o21ai_1 U2 (.A1(n17), .A2(n18), .B1(n16), .Y(carry));
sg13g2_inv_2 U3 (.A(n9), .Y(n13));
sg13g2_o21ai_1 U4 (.A1(n20), .A2(n19), .B1(n14), .Y(n15));
sg13g2_o21ai_1 U5 (.A1(B), .A2(A), .B1(n19), .Y(n18));
sg13g2_nand2_2 U6 (.A(n13), .B(n10), .Y(n12));
sg13g2_inv_2 U7 (.A(n15), .Y(n16));
sg13g2_nand2_2 U8 (.A(n9), .B(cin), .Y(n11));
sg13g2_xnor2_1 U9 (.A(n17), .B(n18), .Y(n9));
sg13g2_nand2_2 U10 (.A(B), .B(A), .Y(n19));
sg13g2_o21ai_1 U11 (.A1(D), .A2(C), .B1(n20), .Y(n17));
sg13g2_nand2_2 U12 (.A(n13), .B(cin), .Y(n14));
sg13g2_nand2_2 U13 (.A(n11), .B(n12), .Y(S));
sg13g2_inv_2 U14 (.A(cin), .Y(n10));
sg13g2_nand2_2 U15 (.A(C), .B(D), .Y(n20));
endmodule

module compressor42_23 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_xnor2_1 U1 (.A(n6), .B(n23), .Y(n5));
sg13g2_inv_2 U2 (.A(n23), .Y(n18));
sg13g2_inv_2 U3 (.A(B), .Y(n10));
sg13g2_nand3_1 U4 (.A(n21), .B(n14), .C(n20), .Y(carry));
sg13g2_nand2_2 U5 (.A(n17), .B(n25), .Y(n6));
sg13g2_nand2_2 U6 (.A(n18), .B(n19), .Y(n20));
sg13g2_inv_2 U7 (.A(C), .Y(n16));
sg13g2_xnor2_1 U8 (.A(n5), .B(cin), .Y(S));
sg13g2_nand2_2 U9 (.A(B), .B(A), .Y(n24));
sg13g2_nand2_2 U10 (.A(n25), .B(n24), .Y(cout));
sg13g2_nand2_2 U11 (.A(n8), .B(cin), .Y(n21));
sg13g2_xnor2_1 U12 (.A(n18), .B(n22), .Y(n8));
sg13g2_nand2_2 U13 (.A(n9), .B(n10), .Y(n11));
sg13g2_nand2_2 U14 (.A(n11), .B(n24), .Y(n23));
sg13g2_inv_2 U15 (.A(A), .Y(n9));
sg13g2_nand2_2 U16 (.A(n15), .B(n16), .Y(n17));
sg13g2_nand2_2 U17 (.A(n12), .B(n13), .Y(n14));
sg13g2_inv_2 U18 (.A(n25), .Y(n12));
sg13g2_inv_2 U19 (.A(n24), .Y(n13));
sg13g2_nand2_2 U20 (.A(n17), .B(n25), .Y(n22));
sg13g2_inv_2 U21 (.A(D), .Y(n15));
sg13g2_inv_2 U22 (.A(n6), .Y(n19));
sg13g2_nand2_2 U23 (.A(D), .B(C), .Y(n25));
endmodule

module compressor42_24 (A, B, C, carry, cin, cout, D, S);
input A, B, C, cin, D;
output carry, cout, S;

sg13g2_nand2_2 U1 (.A(n24), .B(n6), .Y(cout));
sg13g2_inv_2 U2 (.A(n18), .Y(n19));
sg13g2_nand2_2 U3 (.A(n13), .B(n14), .Y(n15));
sg13g2_nand3_1 U4 (.A(n10), .B(n15), .C(n24), .Y(n12));
sg13g2_inv_2 U5 (.A(n22), .Y(n10));
sg13g2_nand3_1 U6 (.A(n17), .B(n1), .C(n20), .Y(carry));
sg13g2_xnor2_1 U7 (.A(n18), .B(cin), .Y(S));
sg13g2_inv_2 U8 (.A(n23), .Y(n5));
sg13g2_inv_2 U9 (.A(n5), .Y(n6));
sg13g2_nand2_2 U10 (.A(B), .B(A), .Y(n23));
sg13g2_nand2_2 U11 (.A(n19), .B(cin), .Y(n20));
sg13g2_o21ai_1 U12 (.A1(A), .A2(B), .B1(n23), .Y(n22));
sg13g2_nand2_2 U13 (.A(D), .B(C), .Y(n24));
sg13g2_nand2_2 U14 (.A(n22), .B(n21), .Y(n11));
sg13g2_nand2_2 U15 (.A(n11), .B(n12), .Y(n18));
sg13g2_nand2_2 U16 (.A(n15), .B(n24), .Y(n21));
sg13g2_inv_2 U17 (.A(D), .Y(n13));
sg13g2_inv_2 U18 (.A(C), .Y(n14));
sg13g2_nand2_2 U19 (.A(n10), .B(n16), .Y(n17));
sg13g2_inv_2 U20 (.A(n21), .Y(n16));
sg13g2_nand2b_1 U21 (.A_N(n24), .B(n5), .Y(n1));
endmodule

module full_adder_0 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n1), .A2(n2), .B1(n3), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n3));
sg13g2_inv_2 U3 (.A(cin), .Y(n2));
sg13g2_xnor2_1 U4 (.A(n1), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n1));
endmodule

module full_adder_1 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(B), .B(A), .Y(n6));
sg13g2_xnor2_1 U5 (.A(cin), .B(n6), .Y(S));
endmodule

module full_adder_2 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(n6), .B(cin), .Y(S));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_o21ai_1 U4 (.A1(n5), .A2(n6), .B1(n4), .Y(cout));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_3 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_inv_2 U1 (.A(n10), .Y(n4));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n8));
sg13g2_inv_2 U3 (.A(cin), .Y(n9));
sg13g2_nand2_2 U4 (.A(n10), .B(cin), .Y(n6));
sg13g2_nand2_2 U5 (.A(n4), .B(n5), .Y(n7));
sg13g2_nand2_2 U6 (.A(n7), .B(n6), .Y(S));
sg13g2_inv_2 U7 (.A(cin), .Y(n5));
sg13g2_o21ai_1 U8 (.A1(n10), .A2(n9), .B1(n8), .Y(cout));
sg13g2_xnor2_1 U9 (.A(B), .B(A), .Y(n10));
endmodule

module full_adder_4 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_inv_2 U1 (.A(n7), .Y(n1));
sg13g2_inv_2 U2 (.A(n1), .Y(n3));
sg13g2_inv_2 U3 (.A(cin), .Y(n4));
sg13g2_xnor2_1 U4 (.A(cin), .B(n9), .Y(S));
sg13g2_nand2_2 U5 (.A(n8), .B(n7), .Y(n9));
sg13g2_nand2_2 U6 (.A(n6), .B(n5), .Y(n8));
sg13g2_nand2_2 U7 (.A(n8), .B(n7), .Y(n10));
sg13g2_inv_2 U8 (.A(A), .Y(n5));
sg13g2_inv_2 U9 (.A(B), .Y(n6));
sg13g2_nand2_2 U10 (.A(A), .B(B), .Y(n7));
sg13g2_o21ai_1 U11 (.A1(n10), .A2(n4), .B1(n3), .Y(cout));
endmodule

module full_adder_5 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(n6), .B(n7), .Y(n9));
sg13g2_nand3_1 U2 (.A(n9), .B(n8), .C(n3), .Y(n5));
sg13g2_nand2_2 U3 (.A(n6), .B(n7), .Y(n1));
sg13g2_inv_2 U4 (.A(B), .Y(n6));
sg13g2_nand2_2 U5 (.A(n2), .B(cin), .Y(n4));
sg13g2_nand2_2 U6 (.A(n1), .B(n8), .Y(n2));
sg13g2_o21ai_1 U7 (.A1(n2), .A2(n3), .B1(n8), .Y(cout));
sg13g2_inv_2 U8 (.A(A), .Y(n7));
sg13g2_nand2_2 U9 (.A(B), .B(A), .Y(n8));
sg13g2_nand2_2 U10 (.A(n5), .B(n4), .Y(S));
sg13g2_inv_2 U11 (.A(cin), .Y(n3));
endmodule

module full_adder_6 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(n2), .B(n4), .Y(net11964));
sg13g2_nand2_2 U2 (.A(n5), .B(A), .Y(n3));
sg13g2_nand2_2 U3 (.A(net11964), .B(net11963), .Y(net12006));
sg13g2_nand2_2 U4 (.A(net11964), .B(net11963), .Y(n1));
sg13g2_inv_2 U5 (.A(B), .Y(n4));
sg13g2_inv_2 U6 (.A(n4), .Y(n5));
sg13g2_inv_2 U7 (.A(A), .Y(n2));
sg13g2_nand2_2 U8 (.A(A), .B(B), .Y(net11963));
sg13g2_nand2_2 U9 (.A(n1), .B(cin), .Y(net10277));
sg13g2_inv_2 U10 (.A(n1), .Y(net10275));
sg13g2_nand2_2 U11 (.A(net10278), .B(net10277), .Y(S));
sg13g2_inv_2 U12 (.A(cin), .Y(net10276));
sg13g2_nand2_2 U13 (.A(net10275), .B(net10276), .Y(net10278));
sg13g2_o21ai_1 U14 (.A1(net10276), .A2(net12006), .B1(n3), .Y(cout));
endmodule

module full_adder_7 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(n6), .B(cin), .Y(S));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_o21ai_1 U4 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_8 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_9 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(n10), .B(cin), .Y(S));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n8));
sg13g2_inv_2 U3 (.A(cin), .Y(n9));
sg13g2_inv_2 U4 (.A(B), .Y(n4));
sg13g2_inv_2 U5 (.A(A), .Y(n5));
sg13g2_o21ai_1 U6 (.A1(n10), .A2(n9), .B1(n8), .Y(cout));
sg13g2_nand2_2 U7 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U8 (.A(n4), .B(n5), .Y(n7));
sg13g2_nand2_2 U9 (.A(n6), .B(n7), .Y(n10));
endmodule

module full_adder_10 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_11 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(n7), .B(n6), .Y(n4));
sg13g2_nand2_2 U2 (.A(n13), .B(n4), .Y(n5));
sg13g2_inv_2 U3 (.A(cin), .Y(n14));
sg13g2_nand2_2 U4 (.A(A), .B(B), .Y(n13));
sg13g2_nand2_2 U5 (.A(n6), .B(n7), .Y(n8));
sg13g2_nand2_2 U6 (.A(n8), .B(n13), .Y(n15));
sg13g2_inv_2 U7 (.A(B), .Y(n6));
sg13g2_inv_2 U8 (.A(A), .Y(n7));
sg13g2_nand2_2 U9 (.A(n5), .B(cin), .Y(n11));
sg13g2_nand2_2 U10 (.A(n9), .B(n10), .Y(n12));
sg13g2_nand2_2 U11 (.A(n11), .B(n12), .Y(S));
sg13g2_inv_2 U12 (.A(n5), .Y(n9));
sg13g2_inv_2 U13 (.A(cin), .Y(n10));
sg13g2_o21ai_1 U14 (.A1(n15), .A2(n14), .B1(n13), .Y(cout));
endmodule

module full_adder_12 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand3_1 U1 (.A(n2), .B(net10321), .C(n5), .Y(n4));
sg13g2_o21ai_1 U2 (.A1(n6), .A2(n2), .B1(n5), .Y(cout));
sg13g2_nand2_2 U3 (.A(n1), .B(cin), .Y(n3));
sg13g2_nand2_2 U4 (.A(n4), .B(n3), .Y(S));
sg13g2_inv_2 U5 (.A(cin), .Y(n2));
sg13g2_inv_2 U6 (.A(net10321), .Y(n6));
sg13g2_inv_2 U7 (.A(B), .Y(net10318));
sg13g2_nand2_2 U8 (.A(net10321), .B(n5), .Y(n1));
sg13g2_nand2_2 U9 (.A(A), .B(B), .Y(n5));
sg13g2_inv_2 U10 (.A(A), .Y(net10319));
sg13g2_nand2_2 U11 (.A(net10318), .B(net10319), .Y(net10321));
endmodule

module full_adder_13 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_inv_2 U1 (.A(B), .Y(n5));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n9));
sg13g2_inv_2 U3 (.A(cin), .Y(n10));
sg13g2_nand2_2 U4 (.A(n7), .B(n8), .Y(n4));
sg13g2_nand2_2 U5 (.A(B), .B(A), .Y(n7));
sg13g2_nand2_2 U6 (.A(n5), .B(n6), .Y(n8));
sg13g2_nand2_2 U7 (.A(n7), .B(n8), .Y(n11));
sg13g2_inv_2 U8 (.A(A), .Y(n6));
sg13g2_o21ai_1 U9 (.A1(n11), .A2(n10), .B1(n9), .Y(cout));
sg13g2_xnor2_1 U10 (.A(cin), .B(n4), .Y(S));
endmodule

module full_adder_14 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand3_1 U1 (.A(n9), .B(n8), .C(n2), .Y(n5));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n10));
sg13g2_inv_2 U3 (.A(A), .Y(n7));
sg13g2_inv_2 U4 (.A(cin), .Y(n2));
sg13g2_inv_2 U5 (.A(B), .Y(n6));
sg13g2_nand2_2 U6 (.A(n11), .B(cin), .Y(n4));
sg13g2_nand2_2 U7 (.A(n5), .B(n4), .Y(S));
sg13g2_nand2_2 U8 (.A(B), .B(A), .Y(n8));
sg13g2_nand2_2 U9 (.A(n7), .B(n6), .Y(n9));
sg13g2_nand2_2 U10 (.A(n9), .B(n8), .Y(n11));
sg13g2_o21ai_1 U11 (.A1(n2), .A2(n11), .B1(n10), .Y(cout));
endmodule

module full_adder_15 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_inv_2 U1 (.A(n6), .Y(n4));
sg13g2_xnor2_1 U2 (.A(cin), .B(n1), .Y(S));
sg13g2_inv_2 U3 (.A(cin), .Y(n11));
sg13g2_nand2_2 U4 (.A(n7), .B(n8), .Y(n1));
sg13g2_inv_2 U5 (.A(B), .Y(n5));
sg13g2_nand2_2 U6 (.A(n4), .B(B), .Y(n10));
sg13g2_inv_2 U7 (.A(A), .Y(n6));
sg13g2_nand2_2 U8 (.A(B), .B(A), .Y(n7));
sg13g2_nand2_2 U9 (.A(n5), .B(n6), .Y(n8));
sg13g2_nand2_2 U10 (.A(n8), .B(n7), .Y(n9));
sg13g2_o21ai_1 U11 (.A1(n9), .A2(n11), .B1(n10), .Y(cout));
endmodule

module full_adder_16 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(net10545), .B(net10546), .Y(n6));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n5));
sg13g2_inv_2 U3 (.A(cin), .Y(n2));
sg13g2_nand2_2 U4 (.A(n6), .B(net10547), .Y(S));
sg13g2_inv_2 U5 (.A(cin), .Y(net10546));
sg13g2_inv_2 U6 (.A(n4), .Y(net10545));
sg13g2_nand2_2 U7 (.A(n4), .B(cin), .Y(net10547));
sg13g2_xnor2_1 U8 (.A(B), .B(A), .Y(n4));
sg13g2_o21ai_1 U9 (.A1(n2), .A2(n4), .B1(n5), .Y(cout));
endmodule

module full_adder_17 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_o21ai_1 U4 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_xnor2_1 U5 (.A(n6), .B(cin), .Y(S));
endmodule

module full_adder_18 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n8));
sg13g2_inv_2 U3 (.A(cin), .Y(n9));
sg13g2_nand2_2 U4 (.A(n4), .B(n5), .Y(n7));
sg13g2_nand2_2 U5 (.A(n6), .B(n7), .Y(n10));
sg13g2_inv_2 U6 (.A(B), .Y(n4));
sg13g2_inv_2 U7 (.A(A), .Y(n5));
sg13g2_xnor2_1 U8 (.A(n10), .B(cin), .Y(S));
sg13g2_o21ai_1 U9 (.A1(n9), .A2(n10), .B1(n8), .Y(cout));
endmodule

module full_adder_19 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n10), .A2(n9), .B1(n8), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n8));
sg13g2_inv_2 U3 (.A(cin), .Y(n9));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U5 (.A(n4), .B(n5), .Y(n7));
sg13g2_nand2_2 U6 (.A(n6), .B(n7), .Y(n10));
sg13g2_inv_2 U7 (.A(B), .Y(n4));
sg13g2_inv_2 U8 (.A(A), .Y(n5));
sg13g2_xnor2_1 U9 (.A(n10), .B(cin), .Y(S));
endmodule

module full_adder_20 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand3_1 U1 (.A(n9), .B(n10), .C(n4), .Y(n6));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n11));
sg13g2_inv_2 U3 (.A(cin), .Y(n12));
sg13g2_nand2_2 U4 (.A(n13), .B(cin), .Y(n5));
sg13g2_nand2_2 U5 (.A(n5), .B(n6), .Y(S));
sg13g2_inv_2 U6 (.A(cin), .Y(n4));
sg13g2_nand2_2 U7 (.A(B), .B(A), .Y(n9));
sg13g2_nand2_2 U8 (.A(n7), .B(n8), .Y(n10));
sg13g2_nand2_2 U9 (.A(n9), .B(n10), .Y(n13));
sg13g2_inv_2 U10 (.A(B), .Y(n7));
sg13g2_inv_2 U11 (.A(A), .Y(n8));
sg13g2_o21ai_1 U12 (.A1(n13), .A2(n12), .B1(n11), .Y(cout));
endmodule

module full_adder_21 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(cin), .B(n2), .Y(S));
sg13g2_nand2_2 U2 (.A(n9), .B(n6), .Y(n2));
sg13g2_nand2_2 U3 (.A(n6), .B(n9), .Y(n10));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n9));
sg13g2_nand2_2 U5 (.A(n4), .B(n5), .Y(n6));
sg13g2_inv_2 U6 (.A(B), .Y(n4));
sg13g2_inv_2 U7 (.A(A), .Y(n5));
sg13g2_inv_2 U8 (.A(n10), .Y(n7));
sg13g2_nand2_2 U9 (.A(n7), .B(cin), .Y(n8));
sg13g2_nand2_2 U10 (.A(n8), .B(n9), .Y(cout));
endmodule

module full_adder_22 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n5), .A2(n6), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_23 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_24 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n7), .A2(n6), .B1(n5), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n5));
sg13g2_inv_2 U3 (.A(cin), .Y(n6));
sg13g2_inv_2 U4 (.A(n6), .Y(n4));
sg13g2_xnor2_1 U5 (.A(n4), .B(n7), .Y(S));
sg13g2_xnor2_1 U6 (.A(B), .B(A), .Y(n7));
endmodule

module full_adder_25 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(n2), .B(n4), .Y(n6));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n7));
sg13g2_o21ai_1 U3 (.A1(n8), .A2(n4), .B1(n7), .Y(cout));
sg13g2_inv_2 U4 (.A(n8), .Y(n2));
sg13g2_nand2_2 U5 (.A(n8), .B(cin), .Y(n5));
sg13g2_nand2_2 U6 (.A(n5), .B(n6), .Y(S));
sg13g2_inv_2 U7 (.A(cin), .Y(n4));
sg13g2_xnor2_1 U8 (.A(B), .B(A), .Y(n8));
endmodule

module full_adder_26 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_27 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_inv_2 U1 (.A(n8), .Y(n2));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n7));
sg13g2_o21ai_1 U3 (.A1(n4), .A2(n8), .B1(n7), .Y(cout));
sg13g2_nand2_2 U4 (.A(n8), .B(cin), .Y(n5));
sg13g2_nand2_2 U5 (.A(n2), .B(n4), .Y(n6));
sg13g2_nand2_2 U6 (.A(n5), .B(n6), .Y(S));
sg13g2_inv_2 U7 (.A(cin), .Y(n4));
sg13g2_xnor2_1 U8 (.A(B), .B(A), .Y(n8));
endmodule

module full_adder_28 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n7), .B1(n5), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n5));
sg13g2_inv_2 U3 (.A(cin), .Y(n6));
sg13g2_xnor2_1 U4 (.A(n7), .B(n4), .Y(S));
sg13g2_xnor2_1 U5 (.A(A), .B(B), .Y(n7));
sg13g2_inv_2 U6 (.A(n6), .Y(n4));
endmodule

module full_adder_29 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_inv_2 U1 (.A(cin), .Y(n3));
sg13g2_nand2_2 U2 (.A(n7), .B(n6), .Y(n9));
sg13g2_inv_2 U3 (.A(A), .Y(n7));
sg13g2_nand2_2 U4 (.A(n10), .B(cin), .Y(n4));
sg13g2_nand2_2 U5 (.A(n2), .B(n3), .Y(n5));
sg13g2_nand2_2 U6 (.A(n5), .B(n4), .Y(S));
sg13g2_inv_2 U7 (.A(n10), .Y(n2));
sg13g2_o21ai_1 U8 (.A1(n10), .A2(n3), .B1(n8), .Y(cout));
sg13g2_nand2_2 U9 (.A(A), .B(B), .Y(n8));
sg13g2_nand2_2 U10 (.A(n8), .B(n9), .Y(n10));
sg13g2_inv_2 U11 (.A(B), .Y(n6));
endmodule

module full_adder_30 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_31 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(n10), .B(cin), .Y(S));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n8));
sg13g2_inv_2 U3 (.A(cin), .Y(n9));
sg13g2_nand2_2 U4 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U5 (.A(n5), .B(n4), .Y(n7));
sg13g2_nand2_2 U6 (.A(n6), .B(n7), .Y(n10));
sg13g2_inv_2 U7 (.A(B), .Y(n4));
sg13g2_inv_2 U8 (.A(A), .Y(n5));
sg13g2_o21ai_1 U9 (.A1(n10), .A2(n9), .B1(n8), .Y(cout));
endmodule

module full_adder_32 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_xnor2_1 U1 (.A(n6), .B(cin), .Y(S));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_o21ai_1 U4 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_33 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n2), .A2(n6), .B1(n5), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n5));
sg13g2_o21ai_1 U3 (.A1(cin), .A2(n6), .B1(n4), .Y(S));
sg13g2_xnor2_1 U4 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U5 (.A(n6), .B(cin), .Y(n4));
sg13g2_inv_2 U6 (.A(cin), .Y(n2));
endmodule

module full_adder_34 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_35 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_36 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_37 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_38 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n7), .A2(n6), .B1(n5), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(n4), .Y(n5));
sg13g2_inv_2 U3 (.A(cin), .Y(n6));
sg13g2_xnor2_1 U4 (.A(n7), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(n4), .B(A), .Y(n7));
sg13g2_buf_2 U6 (.A(B), .X(n4));
endmodule

module full_adder_39 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_40 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_nand2_2 U1 (.A(B), .B(A), .Y(n6));
sg13g2_nand2_2 U2 (.A(B), .B(A), .Y(n8));
sg13g2_inv_2 U3 (.A(cin), .Y(n9));
sg13g2_xnor2_1 U4 (.A(n10), .B(cin), .Y(S));
sg13g2_nand2_2 U5 (.A(n4), .B(n5), .Y(n7));
sg13g2_nand2_2 U6 (.A(n6), .B(n7), .Y(n10));
sg13g2_inv_2 U7 (.A(B), .Y(n4));
sg13g2_inv_2 U8 (.A(A), .Y(n5));
sg13g2_o21ai_1 U9 (.A1(n10), .A2(n9), .B1(n8), .Y(cout));
endmodule

module full_adder_41 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_42 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_43 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module full_adder_44 (A, B, cin, cout, S);
input A, B, cin;
output cout, S;

sg13g2_o21ai_1 U1 (.A1(n6), .A2(n5), .B1(n4), .Y(cout));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(cin), .Y(n5));
sg13g2_xnor2_1 U4 (.A(n6), .B(cin), .Y(S));
sg13g2_xnor2_1 U5 (.A(B), .B(A), .Y(n6));
endmodule

module half_adder_0 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n1), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n1));
sg13g2_xnor2_1 U3 (.A(n2), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n2));
endmodule

module half_adder_1 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_2 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(A), .Y(n6));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n7));
sg13g2_nand2_2 U3 (.A(n6), .B(B), .Y(n4));
sg13g2_inv_2 U4 (.A(B), .Y(n3));
sg13g2_inv_2 U5 (.A(n7), .Y(carry));
sg13g2_nand2_2 U6 (.A(n3), .B(A), .Y(n5));
sg13g2_nand2_2 U7 (.A(n4), .B(n5), .Y(S));
endmodule

module half_adder_3 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_xnor2_1 U1 (.A(n3), .B(B), .Y(S));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U3 (.A(A), .Y(n3));
sg13g2_inv_2 U4 (.A(n4), .Y(carry));
endmodule

module half_adder_4 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(A), .Y(n3));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(n4), .Y(carry));
endmodule

module half_adder_5 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_nand2_2 U1 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U2 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U3 (.A(A), .Y(n3));
sg13g2_inv_2 U4 (.A(n4), .Y(carry));
endmodule

module half_adder_6 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(A), .Y(n6));
sg13g2_nand2_2 U2 (.A(B), .B(n6), .Y(n4));
sg13g2_nand2_2 U3 (.A(n3), .B(A), .Y(n5));
sg13g2_nand2_2 U4 (.A(n4), .B(n5), .Y(S));
sg13g2_inv_2 U5 (.A(B), .Y(n3));
sg13g2_inv_2 U6 (.A(n7), .Y(carry));
sg13g2_nand2_2 U7 (.A(B), .B(A), .Y(n7));
endmodule

module half_adder_7 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_nand2_2 U1 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U2 (.A(n4), .Y(carry));
sg13g2_inv_2 U3 (.A(A), .Y(n3));
sg13g2_xnor2_1 U4 (.A(n3), .B(B), .Y(S));
endmodule

module half_adder_8 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(A), .Y(n3));
sg13g2_xnor2_1 U2 (.A(B), .B(n3), .Y(S));
sg13g2_inv_2 U3 (.A(n4), .Y(carry));
sg13g2_nand2_2 U4 (.A(A), .B(B), .Y(n4));
endmodule

module half_adder_9 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_xnor2_1 U1 (.A(B), .B(n3), .Y(S));
sg13g2_inv_2 U2 (.A(n4), .Y(carry));
sg13g2_nand2_2 U3 (.A(A), .B(B), .Y(n4));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_10 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_11 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_12 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_13 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_14 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_15 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module half_adder_16 (A, B, carry, S);
input A, B;
output carry, S;

sg13g2_inv_2 U1 (.A(n4), .Y(carry));
sg13g2_nand2_2 U2 (.A(A), .B(B), .Y(n4));
sg13g2_xnor2_1 U3 (.A(n3), .B(B), .Y(S));
sg13g2_inv_2 U4 (.A(A), .Y(n3));
endmodule

module partial_product_gen_0 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_nand2_2 U2 (.A(n55), .B(n45), .Y(\pp[10]));
sg13g2_nand2_2 U3 (.A(n53), .B(n43), .Y(n45));
sg13g2_nand2_2 U4 (.A(n58), .B(n41), .Y(\pp[12]));
sg13g2_o21ai_1 U5 (.A1(n7), .A2(n62), .B1(n9), .Y(\pp[8]));
sg13g2_nand2_2 U6 (.A(n53), .B(n2), .Y(n9));
sg13g2_nand2_2 U7 (.A(double), .B(n34), .Y(n8));
sg13g2_inv_2 U8 (.A(n12), .Y(\pp[7]));
sg13g2_inv_2 U9 (.A(n48), .Y(n47));
sg13g2_nor2_2 U10 (.A(n5), .B(n7), .Y(n14));
sg13g2_xnor2_1 U11 (.A(n63), .B(\md[7]), .Y(n7));
sg13g2_inv_2 U12 (.A(n1), .Y(\pp[9]));
sg13g2_a21oi_2 U13 (.A1(n3), .A2(n2), .B1(n4), .Y(n1));
sg13g2_xnor2_1 U14 (.A(n61), .B(\md[6]), .Y(n13));
sg13g2_inv_2 U15 (.A(n17), .Y(\pp[5]));
sg13g2_a21oi_2 U16 (.A1(n18), .A2(n3), .B1(n19), .Y(n17));
sg13g2_nor2_2 U17 (.A(n5), .B(n47), .Y(n19));
sg13g2_xnor2_1 U18 (.A(n63), .B(\md[5]), .Y(n15));
sg13g2_o21ai_1 U19 (.A1(n20), .A2(n62), .B1(n21), .Y(\pp[4]));
sg13g2_nand2_2 U20 (.A(n53), .B(n18), .Y(n21));
sg13g2_xnor2_1 U21 (.A(n60), .B(\md[4]), .Y(n18));
sg13g2_inv_2 U22 (.A(n22), .Y(\pp[3]));
sg13g2_a21oi_2 U23 (.A1(n23), .A2(n3), .B1(n24), .Y(n22));
sg13g2_nor2_2 U24 (.A(n5), .B(n20), .Y(n24));
sg13g2_xnor2_1 U25 (.A(n59), .B(\md[3]), .Y(n20));
sg13g2_o21ai_1 U26 (.A1(n25), .A2(n62), .B1(n26), .Y(\pp[2]));
sg13g2_nand2_2 U27 (.A(n53), .B(n23), .Y(n26));
sg13g2_xnor2_1 U28 (.A(n60), .B(\md[2]), .Y(n23));
sg13g2_inv_2 U29 (.A(n27), .Y(n25));
sg13g2_o21ai_1 U30 (.A1(n28), .A2(n62), .B1(n29), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n53), .B(n27), .Y(n29));
sg13g2_xnor2_1 U32 (.A(n60), .B(\md[1]), .Y(n27));
sg13g2_a21oi_2 U33 (.A1(n3), .A2(n31), .B1(n32), .Y(n30));
sg13g2_nand2_2 U34 (.A(n51), .B(n3), .Y(n52));
sg13g2_nand2_2 U35 (.A(n48), .B(n3), .Y(n49));
sg13g2_a21oi_2 U36 (.A1(n3), .A2(n13), .B1(n14), .Y(n12));
sg13g2_xnor2_1 U37 (.A(n11), .B(\md[15]), .Y(n33));
sg13g2_nor2_2 U38 (.A(n5), .B(n6), .Y(n4));
sg13g2_nand2_2 U39 (.A(n13), .B(n53), .Y(n16));
sg13g2_xnor2_1 U40 (.A(n63), .B(\md[9]), .Y(n6));
sg13g2_nand2_2 U41 (.A(n16), .B(n49), .Y(\pp[6]));
sg13g2_inv_2 U42 (.A(n15), .Y(n48));
sg13g2_xnor2_1 U43 (.A(n60), .B(\md[8]), .Y(n2));
sg13g2_xnor2_1 U44 (.A(negation), .B(\md[13]), .Y(n35));
sg13g2_inv_2 U45 (.A(n30), .Y(\pp[15]));
sg13g2_nand2_2 U46 (.A(n10), .B(n38), .Y(n41));
sg13g2_xnor2_1 U47 (.A(n60), .B(\md[10]), .Y(n43));
sg13g2_inv_2 U48 (.A(n42), .Y(\pp[11]));
sg13g2_a21oi_2 U49 (.A1(n43), .A2(n3), .B1(n44), .Y(n42));
sg13g2_nor2_2 U50 (.A(n5), .B(n40), .Y(n44));
sg13g2_nand2_2 U51 (.A(n53), .B(n31), .Y(n36));
sg13g2_xnor2_1 U52 (.A(n61), .B(\md[14]), .Y(n31));
sg13g2_buf_2 U53 (.A(n64), .X(\pp[16]));
sg13g2_nand2_2 U54 (.A(n56), .B(n34), .Y(n62));
sg13g2_inv_2 U55 (.A(n37), .Y(\pp[13]));
sg13g2_a21oi_2 U56 (.A1(n38), .A2(n3), .B1(n39), .Y(n37));
sg13g2_nor2_2 U57 (.A(n5), .B(n35), .Y(n39));
sg13g2_inv_2 U58 (.A(n10), .Y(n5));
sg13g2_nand2_2 U59 (.A(n52), .B(n36), .Y(\pp[14]));
sg13g2_o21ai_1 U60 (.A1(n28), .A2(n5), .B1(n46), .Y(\pp[0]));
sg13g2_nand2_2 U61 (.A(n56), .B(n59), .Y(n46));
sg13g2_inv_2 U62 (.A(n35), .Y(n51));
sg13g2_xnor2_1 U63 (.A(n61), .B(\md[12]), .Y(n38));
sg13g2_xnor2_1 U64 (.A(n59), .B(\md[0]), .Y(n28));
sg13g2_nand2_2 U65 (.A(n57), .B(n3), .Y(n58));
sg13g2_inv_2 U66 (.A(negation), .Y(n11));
sg13g2_buf_2 U67 (.A(n10), .X(n53));
sg13g2_nand2_2 U68 (.A(n54), .B(n3), .Y(n55));
sg13g2_inv_2 U69 (.A(n6), .Y(n54));
sg13g2_nor2_2 U70 (.A(n64), .B(n56), .Y(n32));
sg13g2_buf_2 U71 (.A(double), .X(n56));
sg13g2_xnor2_1 U72 (.A(n63), .B(\md[11]), .Y(n40));
sg13g2_inv_2 U73 (.A(n40), .Y(n57));
sg13g2_inv_2 U74 (.A(n60), .Y(n59));
sg13g2_nand2_2 U75 (.A(n33), .B(n34), .Y(n64));
sg13g2_buf_2 U76 (.A(n11), .X(n60));
sg13g2_nor2_2 U77 (.A(double), .B(zero), .Y(n10));
sg13g2_buf_2 U78 (.A(n11), .X(n61));
sg13g2_inv_2 U79 (.A(zero), .Y(n34));
sg13g2_buf_2 U80 (.A(negation), .X(n63));
sg13g2_inv_2 U81 (.A(n8), .Y(n3));
endmodule

module partial_product_gen_1 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_xnor2_1 U2 (.A(negation), .B(\md[3]), .Y(n72));
sg13g2_xnor2_1 U3 (.A(n81), .B(\md[2]), .Y(n69));
sg13g2_inv_2 U4 (.A(n75), .Y(\pp[5]));
sg13g2_o21ai_1 U5 (.A1(n85), .A2(n84), .B1(n83), .Y(\pp[8]));
sg13g2_nand2_2 U6 (.A(n82), .B(n90), .Y(n83));
sg13g2_a21oi_2 U7 (.A1(n55), .A2(n89), .B1(n54), .Y(n37));
sg13g2_inv_2 U8 (.A(n80), .Y(\pp[7]));
sg13g2_a21oi_2 U9 (.A1(n79), .A2(n89), .B1(n78), .Y(n80));
sg13g2_nor2_2 U10 (.A(n87), .B(n85), .Y(n78));
sg13g2_xnor2_1 U11 (.A(negation), .B(\md[7]), .Y(n85));
sg13g2_o21ai_1 U12 (.A1(n77), .A2(n84), .B1(n76), .Y(\pp[6]));
sg13g2_nand2_2 U13 (.A(n82), .B(n79), .Y(n76));
sg13g2_xnor2_1 U14 (.A(n81), .B(\md[6]), .Y(n79));
sg13g2_inv_2 U15 (.A(n37), .Y(\pp[13]));
sg13g2_a21oi_2 U16 (.A1(n74), .A2(n89), .B1(n73), .Y(n75));
sg13g2_nor2_2 U17 (.A(n87), .B(n77), .Y(n73));
sg13g2_xnor2_1 U18 (.A(negation), .B(\md[5]), .Y(n77));
sg13g2_o21ai_1 U19 (.A1(n72), .A2(n84), .B1(n71), .Y(\pp[4]));
sg13g2_nand2_2 U20 (.A(n82), .B(n74), .Y(n71));
sg13g2_xnor2_1 U21 (.A(n81), .B(\md[4]), .Y(n74));
sg13g2_inv_2 U22 (.A(n70), .Y(\pp[3]));
sg13g2_a21oi_2 U23 (.A1(n69), .A2(n89), .B1(n68), .Y(n70));
sg13g2_inv_2 U24 (.A(n84), .Y(n89));
sg13g2_nor2_2 U25 (.A(n87), .B(n72), .Y(n68));
sg13g2_nor2_2 U26 (.A(n87), .B(n86), .Y(n88));
sg13g2_nand2_2 U27 (.A(n82), .B(n69), .Y(n66));
sg13g2_xnor2_1 U28 (.A(negation), .B(\md[9]), .Y(n86));
sg13g2_inv_2 U29 (.A(n65), .Y(n67));
sg13g2_o21ai_1 U30 (.A1(n64), .A2(n84), .B1(n63), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n82), .B(n65), .Y(n63));
sg13g2_xnor2_1 U32 (.A(n81), .B(\md[1]), .Y(n65));
sg13g2_inv_2 U33 (.A(n62), .Y(\pp[15]));
sg13g2_a21oi_2 U34 (.A1(n61), .A2(n89), .B1(n60), .Y(n62));
sg13g2_nor2_2 U35 (.A(\pp[16]), .B(double), .Y(n60));
sg13g2_nand2_2 U36 (.A(n59), .B(n58), .Y(\pp[16]));
sg13g2_xnor2_1 U37 (.A(n81), .B(\md[15]), .Y(n59));
sg13g2_o21ai_1 U38 (.A1(n57), .A2(n84), .B1(n56), .Y(\pp[14]));
sg13g2_nand2_2 U39 (.A(n82), .B(n61), .Y(n56));
sg13g2_xnor2_1 U40 (.A(n81), .B(\md[14]), .Y(n61));
sg13g2_inv_2 U41 (.A(negation), .Y(n81));
sg13g2_o21ai_1 U42 (.A1(n67), .A2(n84), .B1(n66), .Y(\pp[2]));
sg13g2_nor2_2 U43 (.A(n87), .B(n57), .Y(n54));
sg13g2_xnor2_1 U44 (.A(negation), .B(\md[13]), .Y(n57));
sg13g2_o21ai_1 U45 (.A1(n53), .A2(n84), .B1(n52), .Y(\pp[12]));
sg13g2_nand2_2 U46 (.A(n82), .B(n55), .Y(n52));
sg13g2_xnor2_1 U47 (.A(n81), .B(\md[12]), .Y(n55));
sg13g2_inv_2 U48 (.A(n51), .Y(\pp[11]));
sg13g2_a21oi_2 U49 (.A1(n50), .A2(n89), .B1(n49), .Y(n51));
sg13g2_nor2_2 U50 (.A(n87), .B(n53), .Y(n49));
sg13g2_xnor2_1 U51 (.A(negation), .B(\md[11]), .Y(n53));
sg13g2_xnor2_1 U52 (.A(n81), .B(\md[8]), .Y(n90));
sg13g2_o21ai_1 U53 (.A1(n86), .A2(n84), .B1(n48), .Y(\pp[10]));
sg13g2_nand2_2 U54 (.A(n82), .B(n50), .Y(n48));
sg13g2_xnor2_1 U55 (.A(n81), .B(\md[10]), .Y(n50));
sg13g2_inv_2 U56 (.A(n91), .Y(\pp[9]));
sg13g2_a21oi_2 U57 (.A1(n90), .A2(n89), .B1(n88), .Y(n91));
sg13g2_nand2_2 U58 (.A(double), .B(n58), .Y(n84));
sg13g2_inv_2 U59 (.A(zero), .Y(n58));
sg13g2_o21ai_1 U60 (.A1(n64), .A2(n87), .B1(n47), .Y(\pp[0]));
sg13g2_nand2_2 U61 (.A(double), .B(negation), .Y(n47));
sg13g2_inv_2 U62 (.A(n82), .Y(n87));
sg13g2_nor2_2 U63 (.A(double), .B(zero), .Y(n82));
sg13g2_xnor2_1 U64 (.A(negation), .B(\md[0]), .Y(n64));
endmodule

module partial_product_gen_2 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_inv_2 U2 (.A(negation), .Y(n88));
sg13g2_xnor2_1 U3 (.A(n88), .B(\md[4]), .Y(n81));
sg13g2_xnor2_1 U4 (.A(negation), .B(\md[13]), .Y(n65));
sg13g2_a21oi_2 U5 (.A1(n96), .A2(n76), .B1(n75), .Y(n77));
sg13g2_nand2_2 U6 (.A(n97), .B(n89), .Y(n90));
sg13g2_a21oi_2 U7 (.A1(n69), .A2(n96), .B1(n68), .Y(n30));
sg13g2_inv_2 U8 (.A(n30), .Y(\pp[15]));
sg13g2_a21oi_2 U9 (.A1(n86), .A2(n96), .B1(n85), .Y(n87));
sg13g2_nor2_2 U10 (.A(n94), .B(n92), .Y(n85));
sg13g2_xnor2_1 U11 (.A(negation), .B(\md[7]), .Y(n92));
sg13g2_o21ai_1 U12 (.A1(n84), .A2(n47), .B1(n83), .Y(\pp[6]));
sg13g2_nand2_2 U13 (.A(n89), .B(n86), .Y(n83));
sg13g2_xnor2_1 U14 (.A(n88), .B(\md[6]), .Y(n86));
sg13g2_o21ai_1 U15 (.A1(n94), .A2(n71), .B1(n54), .Y(\pp[0]));
sg13g2_a21oi_2 U16 (.A1(n81), .A2(n96), .B1(n80), .Y(n82));
sg13g2_nor2_2 U17 (.A(n94), .B(n84), .Y(n80));
sg13g2_xnor2_1 U18 (.A(negation), .B(\md[5]), .Y(n84));
sg13g2_nand2_2 U19 (.A(n67), .B(n66), .Y(\pp[16]));
sg13g2_nand2_2 U20 (.A(n89), .B(n81), .Y(n78));
sg13g2_o21ai_1 U21 (.A1(n60), .A2(n47), .B1(n59), .Y(\pp[12]));
sg13g2_inv_2 U22 (.A(n77), .Y(\pp[3]));
sg13g2_o21ai_1 U23 (.A1(n92), .A2(n47), .B1(n90), .Y(\pp[8]));
sg13g2_nor2_2 U24 (.A(n60), .B(n94), .Y(n56));
sg13g2_inv_2 U25 (.A(n47), .Y(n49));
sg13g2_nand2_2 U26 (.A(n48), .B(n49), .Y(n50));
sg13g2_nand2_2 U27 (.A(n89), .B(n76), .Y(n73));
sg13g2_o21ai_1 U28 (.A1(n74), .A2(n47), .B1(n73), .Y(\pp[2]));
sg13g2_inv_2 U29 (.A(n72), .Y(n74));
sg13g2_o21ai_1 U30 (.A1(n71), .A2(n47), .B1(n70), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n89), .B(n72), .Y(n70));
sg13g2_xnor2_1 U32 (.A(n88), .B(\md[1]), .Y(n72));
sg13g2_inv_2 U33 (.A(n82), .Y(\pp[5]));
sg13g2_xnor2_1 U34 (.A(n88), .B(\md[2]), .Y(n76));
sg13g2_nor2_2 U35 (.A(n94), .B(n79), .Y(n75));
sg13g2_inv_2 U36 (.A(n98), .Y(\pp[9]));
sg13g2_xnor2_1 U37 (.A(n88), .B(\md[15]), .Y(n67));
sg13g2_o21ai_1 U38 (.A1(n65), .A2(n47), .B1(n64), .Y(\pp[14]));
sg13g2_nand2_2 U39 (.A(n89), .B(n69), .Y(n64));
sg13g2_xnor2_1 U40 (.A(n88), .B(\md[14]), .Y(n69));
sg13g2_inv_2 U41 (.A(n93), .Y(n48));
sg13g2_a21oi_2 U42 (.A1(n62), .A2(n96), .B1(n61), .Y(n63));
sg13g2_nor2_2 U43 (.A(n94), .B(n65), .Y(n61));
sg13g2_xnor2_1 U44 (.A(negation), .B(\md[9]), .Y(n93));
sg13g2_nor2_2 U45 (.A(\pp[16]), .B(double), .Y(n68));
sg13g2_nand2_2 U46 (.A(n89), .B(n62), .Y(n59));
sg13g2_xnor2_1 U47 (.A(n88), .B(\md[12]), .Y(n62));
sg13g2_o21ai_1 U48 (.A1(n79), .A2(n47), .B1(n78), .Y(\pp[4]));
sg13g2_a21oi_2 U49 (.A1(n97), .A2(n96), .B1(n95), .Y(n98));
sg13g2_nor2_2 U50 (.A(n94), .B(n93), .Y(n95));
sg13g2_inv_2 U51 (.A(n63), .Y(\pp[13]));
sg13g2_inv_2 U52 (.A(n58), .Y(\pp[11]));
sg13g2_a21oi_2 U53 (.A1(n57), .A2(n96), .B1(n56), .Y(n58));
sg13g2_nand2_2 U54 (.A(n89), .B(n57), .Y(n55));
sg13g2_xnor2_1 U55 (.A(negation), .B(\md[11]), .Y(n60));
sg13g2_xnor2_1 U56 (.A(n88), .B(\md[8]), .Y(n97));
sg13g2_nand2_2 U57 (.A(double), .B(n66), .Y(n47));
sg13g2_nand2_2 U58 (.A(n50), .B(n55), .Y(\pp[10]));
sg13g2_nand2_2 U59 (.A(n88), .B(\md[10]), .Y(n52));
sg13g2_nand2_2 U60 (.A(negation), .B(n51), .Y(n53));
sg13g2_nand2_2 U61 (.A(double), .B(negation), .Y(n54));
sg13g2_nand2_2 U62 (.A(n52), .B(n53), .Y(n57));
sg13g2_inv_2 U63 (.A(\md[10]), .Y(n51));
sg13g2_xnor2_1 U64 (.A(negation), .B(\md[0]), .Y(n71));
sg13g2_xnor2_1 U65 (.A(negation), .B(\md[3]), .Y(n79));
sg13g2_inv_2 U66 (.A(n87), .Y(\pp[7]));
sg13g2_nor2_2 U67 (.A(double), .B(zero), .Y(n89));
sg13g2_inv_2 U68 (.A(zero), .Y(n66));
sg13g2_inv_2 U69 (.A(n91), .Y(n96));
sg13g2_nand2_2 U70 (.A(double), .B(n66), .Y(n91));
sg13g2_inv_2 U71 (.A(n89), .Y(n94));
endmodule

module partial_product_gen_3 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_inv_2 U2 (.A(zero), .Y(n58));
sg13g2_a21oi_2 U3 (.A1(n89), .A2(n61), .B1(n60), .Y(n62));
sg13g2_nor2_2 U4 (.A(\pp[16]), .B(double), .Y(n60));
sg13g2_nand2_2 U5 (.A(n82), .B(n50), .Y(n48));
sg13g2_nand2_2 U6 (.A(n82), .B(n90), .Y(n83));
sg13g2_inv_2 U7 (.A(n91), .Y(\pp[9]));
sg13g2_a21oi_2 U8 (.A1(n89), .A2(n90), .B1(n88), .Y(n91));
sg13g2_a21oi_2 U9 (.A1(n79), .A2(n89), .B1(n78), .Y(n80));
sg13g2_nor2_2 U10 (.A(n87), .B(n85), .Y(n78));
sg13g2_xnor2_1 U11 (.A(negation), .B(\md[7]), .Y(n85));
sg13g2_o21ai_1 U12 (.A1(n77), .A2(n84), .B1(n76), .Y(\pp[6]));
sg13g2_nand2_2 U13 (.A(n82), .B(n79), .Y(n76));
sg13g2_xnor2_1 U14 (.A(n81), .B(\md[6]), .Y(n79));
sg13g2_inv_2 U15 (.A(n75), .Y(\pp[5]));
sg13g2_a21oi_2 U16 (.A1(n74), .A2(n89), .B1(n73), .Y(n75));
sg13g2_inv_2 U17 (.A(n80), .Y(\pp[7]));
sg13g2_inv_2 U18 (.A(n70), .Y(\pp[3]));
sg13g2_o21ai_1 U19 (.A1(n72), .A2(n84), .B1(n71), .Y(\pp[4]));
sg13g2_a21oi_2 U20 (.A1(n89), .A2(n55), .B1(n54), .Y(n37));
sg13g2_inv_2 U21 (.A(n37), .Y(\pp[13]));
sg13g2_nand2_2 U22 (.A(n82), .B(n74), .Y(n71));
sg13g2_a21oi_2 U23 (.A1(n69), .A2(n89), .B1(n68), .Y(n70));
sg13g2_nor2_2 U24 (.A(n87), .B(n72), .Y(n68));
sg13g2_o21ai_1 U25 (.A1(n85), .A2(n84), .B1(n83), .Y(\pp[8]));
sg13g2_inv_2 U26 (.A(negation), .Y(n81));
sg13g2_nand2_2 U27 (.A(n82), .B(n69), .Y(n66));
sg13g2_xnor2_1 U28 (.A(n81), .B(\md[2]), .Y(n69));
sg13g2_inv_2 U29 (.A(n65), .Y(n67));
sg13g2_o21ai_1 U30 (.A1(n64), .A2(n84), .B1(n63), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n82), .B(n65), .Y(n63));
sg13g2_xnor2_1 U32 (.A(n81), .B(\md[1]), .Y(n65));
sg13g2_nand2_2 U33 (.A(n55), .B(n82), .Y(n52));
sg13g2_xnor2_1 U34 (.A(n81), .B(\md[4]), .Y(n74));
sg13g2_xnor2_1 U35 (.A(negation), .B(\md[3]), .Y(n72));
sg13g2_nand2_2 U36 (.A(n59), .B(n58), .Y(\pp[16]));
sg13g2_xnor2_1 U37 (.A(n81), .B(\md[15]), .Y(n59));
sg13g2_o21ai_1 U38 (.A1(n57), .A2(n84), .B1(n56), .Y(\pp[14]));
sg13g2_nand2_2 U39 (.A(n82), .B(n61), .Y(n56));
sg13g2_xnor2_1 U40 (.A(n81), .B(\md[14]), .Y(n61));
sg13g2_inv_2 U41 (.A(n51), .Y(\pp[11]));
sg13g2_o21ai_1 U42 (.A1(n53), .A2(n84), .B1(n52), .Y(\pp[12]));
sg13g2_xnor2_1 U43 (.A(n81), .B(\md[8]), .Y(n90));
sg13g2_nor2_2 U44 (.A(n87), .B(n86), .Y(n88));
sg13g2_a21oi_2 U45 (.A1(n50), .A2(n89), .B1(n49), .Y(n51));
sg13g2_xnor2_1 U46 (.A(n81), .B(\md[10]), .Y(n50));
sg13g2_nor2_2 U47 (.A(n87), .B(n57), .Y(n54));
sg13g2_xnor2_1 U48 (.A(negation), .B(\md[13]), .Y(n57));
sg13g2_nor2_2 U49 (.A(n53), .B(n87), .Y(n49));
sg13g2_xnor2_1 U50 (.A(negation), .B(\md[11]), .Y(n53));
sg13g2_xnor2_1 U51 (.A(n81), .B(\md[12]), .Y(n55));
sg13g2_inv_2 U52 (.A(n62), .Y(\pp[15]));
sg13g2_nor2_2 U53 (.A(n87), .B(n77), .Y(n73));
sg13g2_xnor2_1 U54 (.A(negation), .B(\md[5]), .Y(n77));
sg13g2_o21ai_1 U55 (.A1(n86), .A2(n84), .B1(n48), .Y(\pp[10]));
sg13g2_o21ai_1 U56 (.A1(n67), .A2(n84), .B1(n66), .Y(\pp[2]));
sg13g2_inv_2 U57 (.A(n84), .Y(n89));
sg13g2_xnor2_1 U58 (.A(negation), .B(\md[9]), .Y(n86));
sg13g2_nor2_2 U59 (.A(double), .B(zero), .Y(n82));
sg13g2_o21ai_1 U60 (.A1(n64), .A2(n87), .B1(n47), .Y(\pp[0]));
sg13g2_nand2_2 U61 (.A(double), .B(negation), .Y(n47));
sg13g2_nand2_2 U62 (.A(double), .B(n58), .Y(n84));
sg13g2_inv_2 U63 (.A(n82), .Y(n87));
sg13g2_xnor2_1 U64 (.A(negation), .B(\md[0]), .Y(n64));
endmodule

module partial_product_gen_4 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_inv_2 U2 (.A(n104), .Y(n109));
sg13g2_xnor2_1 U3 (.A(n57), .B(\md[13]), .Y(n78));
sg13g2_a21oi_2 U4 (.A1(n109), .A2(n70), .B1(n69), .Y(n71));
sg13g2_nand2_2 U5 (.A(n80), .B(n79), .Y(\pp[16]));
sg13g2_nand2_2 U6 (.A(n55), .B(n110), .Y(n103));
sg13g2_nand2_2 U7 (.A(n47), .B(n48), .Y(n49));
sg13g2_o21ai_1 U8 (.A1(n11), .A2(n105), .B1(n103), .Y(\pp[8]));
sg13g2_a21oi_2 U9 (.A1(n109), .A2(n100), .B1(n99), .Y(n101));
sg13g2_nor2_2 U10 (.A(n107), .B(n105), .Y(n99));
sg13g2_xnor2_1 U11 (.A(n57), .B(\md[7]), .Y(n105));
sg13g2_o21ai_1 U12 (.A1(n98), .A2(n56), .B1(n97), .Y(\pp[6]));
sg13g2_nand2_2 U13 (.A(n55), .B(n100), .Y(n97));
sg13g2_xnor2_1 U14 (.A(n66), .B(\md[6]), .Y(n100));
sg13g2_inv_2 U15 (.A(n96), .Y(\pp[5]));
sg13g2_a21oi_2 U16 (.A1(n109), .A2(n95), .B1(n94), .Y(n96));
sg13g2_nor2_2 U17 (.A(n107), .B(n98), .Y(n94));
sg13g2_xnor2_1 U18 (.A(n57), .B(\md[5]), .Y(n98));
sg13g2_o21ai_1 U19 (.A1(n93), .A2(n56), .B1(n92), .Y(\pp[4]));
sg13g2_nand2_2 U20 (.A(n55), .B(n95), .Y(n92));
sg13g2_xnor2_1 U21 (.A(n66), .B(\md[4]), .Y(n95));
sg13g2_inv_2 U22 (.A(n91), .Y(\pp[3]));
sg13g2_a21oi_2 U23 (.A1(n109), .A2(n90), .B1(n89), .Y(n91));
sg13g2_nor2_2 U24 (.A(n107), .B(n93), .Y(n89));
sg13g2_xnor2_1 U25 (.A(n57), .B(\md[3]), .Y(n93));
sg13g2_o21ai_1 U26 (.A1(n88), .A2(n11), .B1(n87), .Y(\pp[2]));
sg13g2_nand2_2 U27 (.A(n55), .B(n90), .Y(n87));
sg13g2_xnor2_1 U28 (.A(n66), .B(\md[2]), .Y(n90));
sg13g2_inv_2 U29 (.A(n86), .Y(n88));
sg13g2_o21ai_1 U30 (.A1(n85), .A2(n56), .B1(n84), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n55), .B(n86), .Y(n84));
sg13g2_nor2_2 U32 (.A(n107), .B(n106), .Y(n108));
sg13g2_inv_2 U33 (.A(n58), .Y(n106));
sg13g2_inv_2 U34 (.A(n56), .Y(n48));
sg13g2_inv_2 U35 (.A(n76), .Y(\pp[13]));
sg13g2_inv_2 U36 (.A(n101), .Y(\pp[7]));
sg13g2_inv_2 U37 (.A(n109), .Y(n11));
sg13g2_a21oi_2 U38 (.A1(n82), .A2(n109), .B1(n81), .Y(n83));
sg13g2_xnor2_1 U39 (.A(n65), .B(\md[10]), .Y(n70));
sg13g2_nand2_2 U40 (.A(n82), .B(n55), .Y(n77));
sg13g2_a21oi_2 U41 (.A1(n75), .A2(n109), .B1(n74), .Y(n76));
sg13g2_nor2_2 U42 (.A(n107), .B(n78), .Y(n74));
sg13g2_inv_2 U43 (.A(n83), .Y(\pp[15]));
sg13g2_nor2_2 U44 (.A(\pp[16]), .B(n54), .Y(n81));
sg13g2_nand2_2 U45 (.A(n60), .B(n61), .Y(n80));
sg13g2_nand2_2 U46 (.A(n66), .B(\md[15]), .Y(n60));
sg13g2_nand2_2 U47 (.A(n49), .B(n72), .Y(\pp[12]));
sg13g2_inv_2 U48 (.A(n73), .Y(n47));
sg13g2_nand2_2 U49 (.A(double), .B(n79), .Y(n104));
sg13g2_inv_2 U50 (.A(n111), .Y(\pp[9]));
sg13g2_xnor2_1 U51 (.A(negation), .B(\md[11]), .Y(n73));
sg13g2_xnor2_1 U52 (.A(n66), .B(\md[1]), .Y(n86));
sg13g2_nand2_2 U53 (.A(n62), .B(\md[8]), .Y(n51));
sg13g2_nand2_2 U54 (.A(n64), .B(n50), .Y(n52));
sg13g2_nand2_2 U55 (.A(n51), .B(n52), .Y(n110));
sg13g2_inv_2 U56 (.A(\md[8]), .Y(n50));
sg13g2_a21oi_2 U57 (.A1(n110), .A2(n109), .B1(n108), .Y(n111));
sg13g2_inv_2 U58 (.A(double), .Y(n53));
sg13g2_inv_2 U59 (.A(n53), .Y(n54));
sg13g2_o21ai_1 U60 (.A1(n85), .A2(n107), .B1(n67), .Y(\pp[0]));
sg13g2_nand2_2 U61 (.A(n54), .B(n57), .Y(n67));
sg13g2_nand2_2 U62 (.A(n58), .B(n48), .Y(n63));
sg13g2_nand2_2 U63 (.A(n102), .B(n70), .Y(n68));
sg13g2_xnor2_1 U64 (.A(n57), .B(\md[0]), .Y(n85));
sg13g2_nand2_2 U65 (.A(double), .B(n79), .Y(n56));
sg13g2_xnor2_1 U66 (.A(n65), .B(\md[12]), .Y(n75));
sg13g2_inv_2 U67 (.A(n71), .Y(\pp[11]));
sg13g2_inv_2 U68 (.A(n107), .Y(n55));
sg13g2_inv_2 U69 (.A(negation), .Y(n62));
sg13g2_o21ai_1 U70 (.A1(n78), .A2(n56), .B1(n77), .Y(\pp[14]));
sg13g2_buf_2 U71 (.A(negation), .X(n57));
sg13g2_nand2_2 U72 (.A(n75), .B(n102), .Y(n72));
sg13g2_xnor2_1 U73 (.A(n66), .B(\md[14]), .Y(n82));
sg13g2_inv_2 U74 (.A(n64), .Y(n66));
sg13g2_nor2_2 U75 (.A(n73), .B(n107), .Y(n69));
sg13g2_xnor2_1 U76 (.A(n62), .B(\md[9]), .Y(n58));
sg13g2_nand2_2 U77 (.A(n57), .B(n59), .Y(n61));
sg13g2_inv_2 U78 (.A(\md[15]), .Y(n59));
sg13g2_nand2_2 U79 (.A(n63), .B(n68), .Y(\pp[10]));
sg13g2_inv_2 U80 (.A(n62), .Y(n64));
sg13g2_inv_2 U81 (.A(n64), .Y(n65));
sg13g2_inv_2 U82 (.A(n102), .Y(n107));
sg13g2_nor2_2 U83 (.A(double), .B(zero), .Y(n102));
sg13g2_inv_2 U84 (.A(zero), .Y(n79));
endmodule

module partial_product_gen_5 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_nand2_2 U2 (.A(n48), .B(n89), .Y(n87));
sg13g2_inv_2 U3 (.A(n89), .Y(n51));
sg13g2_inv_2 U4 (.A(n125), .Y(n3));
sg13g2_inv_2 U5 (.A(n3), .Y(\pp[16]));
sg13g2_inv_2 U6 (.A(n92), .Y(n39));
sg13g2_inv_2 U7 (.A(n39), .Y(n47));
sg13g2_inv_2 U8 (.A(zero), .Y(n92));
sg13g2_inv_2 U9 (.A(n113), .Y(n63));
sg13g2_nand2_2 U10 (.A(n116), .B(n113), .Y(n110));
sg13g2_nor2_2 U11 (.A(double), .B(zero), .Y(n48));
sg13g2_o21ai_1 U12 (.A1(n119), .A2(n66), .B1(n117), .Y(\pp[8]));
sg13g2_a21oi_2 U13 (.A1(n108), .A2(n79), .B1(n107), .Y(n109));
sg13g2_nor2_2 U14 (.A(n62), .B(n111), .Y(n107));
sg13g2_inv_2 U15 (.A(\md[14]), .Y(n60));
sg13g2_a21oi_2 U16 (.A1(n85), .A2(n79), .B1(n84), .Y(n86));
sg13g2_inv_2 U17 (.A(\md[0]), .Y(n59));
sg13g2_nor2_2 U18 (.A(n121), .B(n91), .Y(n49));
sg13g2_nand2_2 U19 (.A(n79), .B(n65), .Y(n80));
sg13g2_inv_2 U20 (.A(n49), .Y(n50));
sg13g2_o21ai_1 U21 (.A1(n51), .A2(n52), .B1(n50), .Y(\pp[13]));
sg13g2_inv_2 U22 (.A(n79), .Y(n52));
sg13g2_nor2_2 U23 (.A(n62), .B(n106), .Y(n102));
sg13g2_inv_2 U24 (.A(n65), .Y(n106));
sg13g2_inv_2 U25 (.A(n79), .Y(n77));
sg13g2_nand2_2 U26 (.A(n93), .B(n47), .Y(n125));
sg13g2_nand2_2 U27 (.A(n61), .B(n103), .Y(n100));
sg13g2_inv_2 U28 (.A(n114), .Y(\pp[7]));
sg13g2_inv_2 U29 (.A(n99), .Y(n101));
sg13g2_o21ai_1 U30 (.A1(n66), .A2(n98), .B1(n97), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n61), .B(n99), .Y(n97));
sg13g2_xnor2_1 U32 (.A(n115), .B(\md[1]), .Y(n99));
sg13g2_nor2_2 U33 (.A(n125), .B(n75), .Y(n94));
sg13g2_nand2_2 U34 (.A(n61), .B(n123), .Y(n117));
sg13g2_xnor2_1 U35 (.A(n115), .B(\md[12]), .Y(n89));
sg13g2_nand2_2 U36 (.A(n55), .B(n56), .Y(n58));
sg13g2_inv_2 U37 (.A(n55), .Y(n53));
sg13g2_inv_2 U38 (.A(negation), .Y(n55));
sg13g2_nand2_2 U39 (.A(n53), .B(\md[7]), .Y(n73));
sg13g2_inv_2 U40 (.A(n53), .Y(n71));
sg13g2_xnor2_1 U41 (.A(n81), .B(n60), .Y(n95));
sg13g2_inv_2 U42 (.A(n115), .Y(n81));
sg13g2_nor2_2 U43 (.A(n119), .B(n62), .Y(n112));
sg13g2_o21ai_1 U44 (.A1(n98), .A2(n62), .B1(n82), .Y(\pp[0]));
sg13g2_xnor2_1 U45 (.A(n115), .B(n59), .Y(n98));
sg13g2_xnor2_1 U46 (.A(n115), .B(\md[4]), .Y(n108));
sg13g2_inv_2 U47 (.A(n124), .Y(\pp[9]));
sg13g2_a21oi_2 U48 (.A1(n123), .A2(n79), .B1(n122), .Y(n124));
sg13g2_nor2_2 U49 (.A(n63), .B(n77), .Y(n64));
sg13g2_inv_2 U50 (.A(\md[8]), .Y(n54));
sg13g2_xnor2_1 U51 (.A(n53), .B(n54), .Y(n123));
sg13g2_inv_2 U52 (.A(n62), .Y(n61));
sg13g2_nor2_2 U53 (.A(n76), .B(n77), .Y(n78));
sg13g2_nand2_2 U54 (.A(n116), .B(n85), .Y(n83));
sg13g2_inv_2 U55 (.A(n104), .Y(\pp[3]));
sg13g2_xnor2_1 U56 (.A(n115), .B(\md[6]), .Y(n113));
sg13g2_nand2_2 U57 (.A(n61), .B(n95), .Y(n90));
sg13g2_inv_2 U58 (.A(n86), .Y(\pp[11]));
sg13g2_nand2_2 U59 (.A(negation), .B(\md[9]), .Y(n57));
sg13g2_nand2_2 U60 (.A(n57), .B(n58), .Y(n120));
sg13g2_nand2_2 U61 (.A(n75), .B(negation), .Y(n82));
sg13g2_inv_2 U62 (.A(\md[9]), .Y(n56));
sg13g2_o21ai_1 U63 (.A1(n120), .A2(n77), .B1(n83), .Y(\pp[10]));
sg13g2_inv_2 U64 (.A(n118), .Y(n79));
sg13g2_nor2_2 U65 (.A(n121), .B(n88), .Y(n84));
sg13g2_nand2_2 U66 (.A(n61), .B(n108), .Y(n105));
sg13g2_a21oi_2 U67 (.A1(n95), .A2(n79), .B1(n94), .Y(n96));
sg13g2_nand2_2 U68 (.A(n105), .B(n80), .Y(\pp[4]));
sg13g2_o21ai_1 U69 (.A1(n77), .A2(n88), .B1(n87), .Y(\pp[12]));
sg13g2_o21ai_1 U70 (.A1(n91), .A2(n66), .B1(n90), .Y(\pp[14]));
sg13g2_xnor2_1 U71 (.A(negation), .B(\md[13]), .Y(n91));
sg13g2_inv_2 U72 (.A(n48), .Y(n62));
sg13g2_nor2_2 U73 (.A(n102), .B(n78), .Y(n104));
sg13g2_nor2_2 U74 (.A(n112), .B(n64), .Y(n114));
sg13g2_xnor2_1 U75 (.A(n115), .B(\md[3]), .Y(n65));
sg13g2_nor2_2 U76 (.A(n121), .B(n120), .Y(n122));
sg13g2_buf_2 U77 (.A(n118), .X(n66));
sg13g2_xnor2_1 U78 (.A(n115), .B(\md[15]), .Y(n93));
sg13g2_inv_2 U79 (.A(n103), .Y(n76));
sg13g2_nand2_2 U80 (.A(n115), .B(\md[10]), .Y(n69));
sg13g2_nand2_2 U81 (.A(n81), .B(n68), .Y(n70));
sg13g2_nand2_2 U82 (.A(n69), .B(n70), .Y(n85));
sg13g2_inv_2 U83 (.A(\md[10]), .Y(n68));
sg13g2_xnor2_1 U84 (.A(n115), .B(\md[2]), .Y(n103));
sg13g2_nand2_2 U85 (.A(n71), .B(n72), .Y(n74));
sg13g2_nand2_2 U86 (.A(n73), .B(n74), .Y(n119));
sg13g2_inv_2 U87 (.A(\md[7]), .Y(n72));
sg13g2_inv_2 U88 (.A(n109), .Y(\pp[5]));
sg13g2_o21ai_1 U89 (.A1(n111), .A2(n66), .B1(n110), .Y(\pp[6]));
sg13g2_buf_2 U90 (.A(double), .X(n75));
sg13g2_inv_2 U91 (.A(n96), .Y(\pp[15]));
sg13g2_xnor2_1 U92 (.A(negation), .B(\md[11]), .Y(n88));
sg13g2_xnor2_1 U93 (.A(n81), .B(\md[5]), .Y(n111));
sg13g2_o21ai_1 U94 (.A1(n101), .A2(n66), .B1(n100), .Y(\pp[2]));
sg13g2_inv_2 U95 (.A(negation), .Y(n115));
sg13g2_nand2_2 U96 (.A(n92), .B(double), .Y(n118));
sg13g2_inv_2 U97 (.A(n116), .Y(n121));
sg13g2_nor2_2 U98 (.A(double), .B(zero), .Y(n116));
endmodule

module partial_product_gen_6 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_inv_2 U2 (.A(n116), .Y(n25));
sg13g2_nand2_2 U3 (.A(negation), .B(n50), .Y(n52));
sg13g2_nand2_2 U4 (.A(negation), .B(n47), .Y(n49));
sg13g2_nand2_2 U5 (.A(n73), .B(n101), .Y(n98));
sg13g2_inv_2 U6 (.A(n72), .Y(n73));
sg13g2_inv_2 U7 (.A(n89), .Y(n54));
sg13g2_inv_2 U8 (.A(n77), .Y(n58));
sg13g2_xnor2_1 U9 (.A(n108), .B(\md[10]), .Y(n77));
sg13g2_o21ai_1 U10 (.A1(n104), .A2(n69), .B1(n103), .Y(\pp[6]));
sg13g2_inv_2 U11 (.A(n60), .Y(n93));
sg13g2_a21oi_2 U12 (.A1(n116), .A2(n101), .B1(n100), .Y(n102));
sg13g2_nor2_2 U13 (.A(n71), .B(\pp[16]), .Y(n88));
sg13g2_nand2_2 U14 (.A(n71), .B(n68), .Y(n74));
sg13g2_inv_2 U15 (.A(n70), .Y(n71));
sg13g2_nor2_2 U16 (.A(n114), .B(n113), .Y(n115));
sg13g2_a21oi_2 U17 (.A1(n116), .A2(n96), .B1(n95), .Y(n97));
sg13g2_nor2_2 U18 (.A(n114), .B(n99), .Y(n95));
sg13g2_inv_2 U19 (.A(zero), .Y(n86));
sg13g2_inv_2 U20 (.A(n111), .Y(n116));
sg13g2_inv_2 U21 (.A(n116), .Y(n53));
sg13g2_inv_2 U22 (.A(n97), .Y(\pp[3]));
sg13g2_inv_2 U23 (.A(negation), .Y(n108));
sg13g2_xnor2_1 U24 (.A(negation), .B(\md[5]), .Y(n104));
sg13g2_nand2_2 U25 (.A(n108), .B(\md[15]), .Y(n48));
sg13g2_nand2_2 U26 (.A(n48), .B(n49), .Y(n87));
sg13g2_inv_2 U27 (.A(\md[15]), .Y(n47));
sg13g2_xnor2_1 U28 (.A(n108), .B(\md[12]), .Y(n82));
sg13g2_nor2_2 U29 (.A(n114), .B(n104), .Y(n100));
sg13g2_o21ai_1 U30 (.A1(n92), .A2(n69), .B1(n91), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(n73), .B(n93), .Y(n91));
sg13g2_inv_2 U32 (.A(n73), .Y(n114));
sg13g2_inv_2 U33 (.A(n85), .Y(n65));
sg13g2_o21ai_1 U34 (.A1(n80), .A2(n53), .B1(n79), .Y(\pp[12]));
sg13g2_nand2_2 U35 (.A(n108), .B(\md[8]), .Y(n51));
sg13g2_nand2_2 U36 (.A(n51), .B(n52), .Y(n117));
sg13g2_inv_2 U37 (.A(\md[8]), .Y(n50));
sg13g2_nor2_2 U38 (.A(n114), .B(n112), .Y(n105));
sg13g2_nand2_2 U39 (.A(n73), .B(n96), .Y(n94));
sg13g2_inv_2 U40 (.A(n82), .Y(n56));
sg13g2_a21oi_2 U41 (.A1(n106), .A2(n116), .B1(n105), .Y(n107));
sg13g2_inv_2 U42 (.A(n102), .Y(\pp[5]));
sg13g2_nor2_2 U43 (.A(n25), .B(n54), .Y(n55));
sg13g2_nor2_2 U44 (.A(n55), .B(n88), .Y(n90));
sg13g2_xnor2_1 U45 (.A(n108), .B(\md[2]), .Y(n96));
sg13g2_nand2_2 U46 (.A(n73), .B(n82), .Y(n79));
sg13g2_nor2_2 U47 (.A(n56), .B(n25), .Y(n57));
sg13g2_nor2_2 U48 (.A(n81), .B(n57), .Y(n83));
sg13g2_inv_2 U49 (.A(n83), .Y(\pp[13]));
sg13g2_o21ai_1 U50 (.A1(n69), .A2(n113), .B1(n75), .Y(\pp[10]));
sg13g2_nor2_2 U51 (.A(n58), .B(n53), .Y(n59));
sg13g2_nor2_2 U52 (.A(n59), .B(n76), .Y(n78));
sg13g2_nor2_2 U53 (.A(n114), .B(n80), .Y(n76));
sg13g2_nand2_2 U54 (.A(n73), .B(n77), .Y(n75));
sg13g2_inv_2 U55 (.A(n90), .Y(\pp[15]));
sg13g2_inv_2 U56 (.A(n118), .Y(\pp[9]));
sg13g2_xnor2_1 U57 (.A(negation), .B(\md[11]), .Y(n80));
sg13g2_a21oi_2 U58 (.A1(n117), .A2(n116), .B1(n115), .Y(n118));
sg13g2_xnor2_1 U59 (.A(n61), .B(\md[1]), .Y(n60));
sg13g2_o21ai_1 U60 (.A1(n92), .A2(n114), .B1(n74), .Y(\pp[0]));
sg13g2_inv_2 U61 (.A(n108), .Y(n61));
sg13g2_nor2_2 U62 (.A(n114), .B(n85), .Y(n81));
sg13g2_xnor2_1 U63 (.A(n108), .B(\md[4]), .Y(n101));
sg13g2_xnor2_1 U64 (.A(n61), .B(\md[0]), .Y(n92));
sg13g2_xnor2_1 U65 (.A(n68), .B(\md[7]), .Y(n112));
sg13g2_o21ai_1 U66 (.A1(n99), .A2(n69), .B1(n98), .Y(\pp[4]));
sg13g2_xnor2_1 U67 (.A(n61), .B(\md[3]), .Y(n99));
sg13g2_nand2_2 U68 (.A(n73), .B(n106), .Y(n103));
sg13g2_inv_2 U69 (.A(n109), .Y(n72));
sg13g2_o21ai_1 U70 (.A1(n60), .A2(n69), .B1(n94), .Y(\pp[2]));
sg13g2_inv_2 U71 (.A(n78), .Y(\pp[11]));
sg13g2_nand2_2 U72 (.A(n86), .B(n87), .Y(\pp[16]));
sg13g2_nand2_2 U73 (.A(n68), .B(\md[13]), .Y(n63));
sg13g2_nand2_2 U74 (.A(n108), .B(n62), .Y(n64));
sg13g2_nand2_2 U75 (.A(n63), .B(n64), .Y(n85));
sg13g2_inv_2 U76 (.A(\md[13]), .Y(n62));
sg13g2_o21ai_1 U77 (.A1(n112), .A2(n69), .B1(n110), .Y(\pp[8]));
sg13g2_nand2_2 U78 (.A(n73), .B(n117), .Y(n110));
sg13g2_inv_2 U79 (.A(n107), .Y(\pp[7]));
sg13g2_xnor2_1 U80 (.A(n108), .B(\md[14]), .Y(n89));
sg13g2_nand2_2 U81 (.A(n65), .B(n66), .Y(n67));
sg13g2_nand2_2 U82 (.A(n67), .B(n84), .Y(\pp[14]));
sg13g2_inv_2 U83 (.A(n69), .Y(n66));
sg13g2_nand2_2 U84 (.A(n73), .B(n89), .Y(n84));
sg13g2_xnor2_1 U85 (.A(n108), .B(\md[6]), .Y(n106));
sg13g2_buf_2 U86 (.A(negation), .X(n68));
sg13g2_xnor2_1 U87 (.A(negation), .B(\md[9]), .Y(n113));
sg13g2_buf_2 U88 (.A(n111), .X(n69));
sg13g2_inv_2 U89 (.A(double), .Y(n70));
sg13g2_nand2_2 U90 (.A(n86), .B(double), .Y(n111));
sg13g2_nor2_2 U91 (.A(double), .B(zero), .Y(n109));
endmodule

module partial_product_gen_7 (\md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16], double, negation, zero);
input \md[0], \md[1], \md[2], \md[3], \md[4], \md[5], \md[6], \md[7], \md[8], \md[9], \md[10], \md[11], \md[12], \md[13], \md[14], \md[15], double, negation, zero;
output \pp[0], \pp[1], \pp[2], \pp[3], \pp[4], \pp[5], \pp[6], \pp[7], \pp[8], \pp[9], \pp[10], \pp[11], \pp[12], \pp[13], \pp[14], \pp[15], \pp[16];

sg13g2_o21ai_1 U2 (.A1(n98), .A2(n8), .B1(n97), .Y(\pp[8]));
sg13g2_a21oi_2 U3 (.A1(n58), .A2(n101), .B1(n100), .Y(n102));
sg13g2_o21ai_1 U4 (.A1(n99), .A2(n8), .B1(n45), .Y(\pp[10]));
sg13g2_nand2_2 U5 (.A(n3), .B(n64), .Y(n66));
sg13g2_inv_2 U6 (.A(n96), .Y(\pp[7]));
sg13g2_inv_2 U7 (.A(n56), .Y(n3));
sg13g2_a21oi_2 U8 (.A1(n13), .A2(n58), .B1(n95), .Y(n96));
sg13g2_o21ai_1 U9 (.A1(n69), .A2(n8), .B1(n68), .Y(\pp[12]));
sg13g2_nand2_2 U10 (.A(n62), .B(n58), .Y(n63));
sg13g2_inv_2 U11 (.A(n74), .Y(n62));
sg13g2_o21ai_1 U12 (.A1(n94), .A2(n8), .B1(n93), .Y(\pp[6]));
sg13g2_nand2_2 U13 (.A(net10722), .B(n13), .Y(n93));
sg13g2_nand2_2 U14 (.A(n60), .B(n58), .Y(n61));
sg13g2_inv_2 U15 (.A(n92), .Y(\pp[5]));
sg13g2_a21oi_2 U16 (.A1(n91), .A2(n58), .B1(n90), .Y(n92));
sg13g2_nor2_2 U17 (.A(n5), .B(n94), .Y(n90));
sg13g2_xnor2_1 U18 (.A(n57), .B(\md[5]), .Y(n94));
sg13g2_nor2_2 U19 (.A(n5), .B(n99), .Y(n100));
sg13g2_nor2_2 U20 (.A(n103), .B(n47), .Y(n77));
sg13g2_inv_2 U21 (.A(n79), .Y(\pp[15]));
sg13g2_inv_2 U22 (.A(n87), .Y(\pp[3]));
sg13g2_a21oi_2 U23 (.A1(n86), .A2(n58), .B1(n85), .Y(n87));
sg13g2_nor2_2 U24 (.A(n5), .B(n89), .Y(n85));
sg13g2_inv_2 U25 (.A(n102), .Y(\pp[9]));
sg13g2_o21ai_1 U26 (.A1(n84), .A2(n48), .B1(n83), .Y(\pp[2]));
sg13g2_nand2_2 U27 (.A(net10722), .B(n86), .Y(n83));
sg13g2_xnor2_1 U28 (.A(n11), .B(\md[2]), .Y(n86));
sg13g2_inv_2 U29 (.A(n82), .Y(n84));
sg13g2_o21ai_1 U30 (.A1(n81), .A2(n48), .B1(n80), .Y(\pp[1]));
sg13g2_nand2_2 U31 (.A(net10722), .B(n82), .Y(n80));
sg13g2_xnor2_1 U32 (.A(n11), .B(\md[1]), .Y(n82));
sg13g2_nand2_2 U33 (.A(net10722), .B(n53), .Y(n45));
sg13g2_xnor2_1 U34 (.A(n57), .B(\md[9]), .Y(n99));
sg13g2_xnor2_1 U35 (.A(n57), .B(\md[3]), .Y(n89));
sg13g2_nor2_2 U36 (.A(n54), .B(n8), .Y(n52));
sg13g2_inv_2 U37 (.A(double), .Y(n43));
sg13g2_inv_2 U38 (.A(n43), .Y(n47));
sg13g2_xnor2_1 U39 (.A(n57), .B(\md[10]), .Y(n54));
sg13g2_inv_2 U40 (.A(n58), .Y(n48));
sg13g2_inv_2 U41 (.A(n49), .Y(n50));
sg13g2_nand2_2 U42 (.A(net10722), .B(n78), .Y(n73));
sg13g2_nor2_2 U43 (.A(n69), .B(n5), .Y(n44));
sg13g2_nand2_2 U44 (.A(n76), .B(n50), .Y(n103));
sg13g2_inv_2 U45 (.A(n42), .Y(\pp[11]));
sg13g2_inv_2 U46 (.A(n75), .Y(n49));
sg13g2_xnor2_1 U47 (.A(n57), .B(\md[13]), .Y(n74));
sg13g2_nor2_2 U48 (.A(n52), .B(n44), .Y(n42));
sg13g2_xnor2_1 U49 (.A(n11), .B(\md[15]), .Y(n76));
sg13g2_inv_2 U50 (.A(n54), .Y(n53));
sg13g2_xnor2_1 U51 (.A(n11), .B(\md[8]), .Y(n101));
sg13g2_nand2_2 U52 (.A(n101), .B(net10722), .Y(n97));
sg13g2_inv_2 U53 (.A(n55), .Y(n13));
sg13g2_xnor2_1 U54 (.A(n56), .B(\md[4]), .Y(n91));
sg13g2_a21oi_2 U55 (.A1(n58), .A2(n78), .B1(n77), .Y(n79));
sg13g2_inv_2 U56 (.A(n8), .Y(n58));
sg13g2_nor2_2 U57 (.A(double), .B(zero), .Y(n51));
sg13g2_nor2_2 U58 (.A(double), .B(zero), .Y(n10));
sg13g2_nor2_2 U59 (.A(n5), .B(n98), .Y(n95));
sg13g2_o21ai_1 U60 (.A1(n81), .A2(n5), .B1(n67), .Y(\pp[0]));
sg13g2_nand2_2 U61 (.A(n47), .B(net9683), .Y(n67));
sg13g2_xnor2_1 U62 (.A(n57), .B(\md[6]), .Y(n55));
sg13g2_inv_2 U63 (.A(n56), .Y(n57));
sg13g2_xnor2_1 U64 (.A(n57), .B(\md[0]), .Y(n81));
sg13g2_inv_2 U65 (.A(negation), .Y(n56));
sg13g2_inv_2 U66 (.A(n51), .Y(n5));
sg13g2_nand2_2 U67 (.A(n76), .B(n50), .Y(\pp[16]));
sg13g2_nand2_2 U68 (.A(n11), .B(\md[12]), .Y(n65));
sg13g2_nand2_2 U69 (.A(net10722), .B(n71), .Y(n68));
sg13g2_nand2_2 U70 (.A(n61), .B(n88), .Y(\pp[4]));
sg13g2_inv_2 U71 (.A(n89), .Y(n60));
sg13g2_inv_2 U72 (.A(n72), .Y(\pp[13]));
sg13g2_a21oi_2 U73 (.A1(n71), .A2(n58), .B1(n70), .Y(n72));
sg13g2_nand2_2 U74 (.A(net10722), .B(n91), .Y(n88));
sg13g2_nor2_2 U75 (.A(n5), .B(n74), .Y(n70));
sg13g2_xnor2_1 U76 (.A(n57), .B(\md[7]), .Y(n98));
sg13g2_xnor2_1 U77 (.A(n57), .B(\md[11]), .Y(n69));
sg13g2_inv_2 U78 (.A(zero), .Y(n75));
sg13g2_nand2_2 U79 (.A(n63), .B(n73), .Y(\pp[14]));
sg13g2_xnor2_1 U80 (.A(n11), .B(\md[14]), .Y(n78));
sg13g2_buf_2 U81 (.A(n10), .X(net10722));
sg13g2_inv_2 U82 (.A(negation), .Y(n11));
sg13g2_nand2_2 U83 (.A(n65), .B(n66), .Y(n71));
sg13g2_inv_2 U84 (.A(n11), .Y(net9683));
sg13g2_inv_2 U85 (.A(\md[12]), .Y(n64));
sg13g2_nand2_2 U86 (.A(double), .B(n75), .Y(n8));
endmodule

