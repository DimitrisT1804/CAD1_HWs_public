// Generated netlist by CADI API on Date: 2025-10-09 17:33:06 //

module c499 (N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755);
input N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;

sg13g2_xor2_1 U186 (.A(N125), .B(n154), .X(N755));
sg13g2_nor2_1 U187 (.A(n155), .B(n156), .Y(n154));
sg13g2_xor2_1 U188 (.A(N121), .B(n157), .X(N754));
sg13g2_nor2_1 U189 (.A(n158), .B(n156), .Y(n157));
sg13g2_xor2_1 U190 (.A(N117), .B(n159), .X(N753));
sg13g2_nor2_1 U191 (.A(n160), .B(n156), .Y(n159));
sg13g2_xor2_1 U192 (.A(N113), .B(n161), .X(N752));
sg13g2_nor2_1 U193 (.A(n162), .B(n156), .Y(n161));
sg13g2_nand4_1 U194 (.A(n163), .B(n164), .C(n165), .D(n166), .Y(n156));
sg13g2_xor2_1 U195 (.A(N109), .B(n167), .X(N751));
sg13g2_nor2_1 U196 (.A(n155), .B(n168), .Y(n167));
sg13g2_xor2_1 U197 (.A(N105), .B(n169), .X(N750));
sg13g2_nor2_1 U198 (.A(n158), .B(n168), .Y(n169));
sg13g2_xor2_1 U199 (.A(N101), .B(n170), .X(N749));
sg13g2_nor2_1 U200 (.A(n160), .B(n168), .Y(n170));
sg13g2_xor2_1 U201 (.A(N97), .B(n171), .X(N748));
sg13g2_nor2_1 U202 (.A(n162), .B(n168), .Y(n171));
sg13g2_nand4_1 U203 (.A(n172), .B(n166), .C(n173), .D(n174), .Y(n168));
sg13g2_nor2_1 U204 (.A(n175), .B(n176), .Y(n174));
sg13g2_xor2_1 U205 (.A(N93), .B(n177), .X(N747));
sg13g2_nor2_1 U206 (.A(n155), .B(n178), .Y(n177));
sg13g2_xor2_1 U207 (.A(N89), .B(n179), .X(N746));
sg13g2_nor2_1 U208 (.A(n158), .B(n178), .Y(n179));
sg13g2_xor2_1 U209 (.A(N85), .B(n180), .X(N745));
sg13g2_nor2_1 U210 (.A(n160), .B(n178), .Y(n180));
sg13g2_xor2_1 U211 (.A(N81), .B(n181), .X(N744));
sg13g2_nor2_1 U212 (.A(n162), .B(n178), .Y(n181));
sg13g2_nand4_1 U213 (.A(n176), .B(n166), .C(n175), .D(n182), .Y(n178));
sg13g2_nor2_1 U214 (.A(n173), .B(n172), .Y(n182));
sg13g2_xor2_1 U215 (.A(N77), .B(n183), .X(N743));
sg13g2_nor2_1 U216 (.A(n155), .B(n184), .Y(n183));
sg13g2_xor2_1 U217 (.A(N73), .B(n185), .X(N742));
sg13g2_nor2_1 U218 (.A(n158), .B(n184), .Y(n185));
sg13g2_xor2_1 U219 (.A(N69), .B(n186), .X(N741));
sg13g2_nor2_1 U220 (.A(n160), .B(n184), .Y(n186));
sg13g2_xor2_1 U221 (.A(N65), .B(n187), .X(N740));
sg13g2_nor2_1 U222 (.A(n162), .B(n184), .Y(n187));
sg13g2_nand4_1 U223 (.A(n188), .B(n189), .C(n190), .D(n166), .Y(n184));
sg13g2_nand2_1 U224 (.A(n191), .B(n192), .Y(n166));
sg13g2_or3_1 U225 (.A(n193), .B(n194), .C(n195), .X(n192));
sg13g2_or3_1 U226 (.A(n196), .B(n197), .C(n198), .X(n191));
sg13g2_xor2_1 U227 (.A(N61), .B(n199), .X(N739));
sg13g2_nor2_1 U228 (.A(n190), .B(n200), .Y(n199));
sg13g2_xor2_1 U229 (.A(N57), .B(n201), .X(N738));
sg13g2_nor2_1 U230 (.A(n165), .B(n200), .Y(n201));
sg13g2_xor2_1 U231 (.A(N53), .B(n202), .X(N737));
sg13g2_nor2_1 U232 (.A(n188), .B(n200), .Y(n202));
sg13g2_xor2_1 U233 (.A(N49), .B(n203), .X(N736));
sg13g2_nor2_1 U234 (.A(n163), .B(n200), .Y(n203));
sg13g2_nand4_1 U235 (.A(n158), .B(n196), .C(n162), .D(n204), .Y(n200));
sg13g2_nor2_1 U236 (.A(n160), .B(n155), .Y(n196));
sg13g2_xor2_1 U237 (.A(N45), .B(n205), .X(N735));
sg13g2_nor2_1 U238 (.A(n190), .B(n206), .Y(n205));
sg13g2_xor2_1 U239 (.A(N41), .B(n207), .X(N734));
sg13g2_nor2_1 U240 (.A(n165), .B(n206), .Y(n207));
sg13g2_xor2_1 U241 (.A(N37), .B(n208), .X(N733));
sg13g2_nor2_1 U242 (.A(n188), .B(n206), .Y(n208));
sg13g2_xor2_1 U243 (.A(N33), .B(n209), .X(N732));
sg13g2_nor2_1 U244 (.A(n163), .B(n206), .Y(n209));
sg13g2_nand4_1 U245 (.A(n198), .B(n204), .C(n194), .D(n210), .Y(n206));
sg13g2_nor2_1 U246 (.A(n195), .B(n197), .Y(n210));
sg13g2_xor2_1 U247 (.A(N29), .B(n211), .X(N731));
sg13g2_nor2_1 U248 (.A(n190), .B(n212), .Y(n211));
sg13g2_xor2_1 U249 (.A(N25), .B(n213), .X(N730));
sg13g2_nor2_1 U250 (.A(n165), .B(n212), .Y(n213));
sg13g2_xor2_1 U251 (.A(N21), .B(n214), .X(N729));
sg13g2_nor2_1 U252 (.A(n188), .B(n212), .Y(n214));
sg13g2_xor2_1 U253 (.A(N17), .B(n215), .X(N728));
sg13g2_nor2_1 U254 (.A(n163), .B(n212), .Y(n215));
sg13g2_nand4_1 U255 (.A(n197), .B(n204), .C(n195), .D(n216), .Y(n212));
sg13g2_nor2_1 U256 (.A(n198), .B(n194), .Y(n216));
sg13g2_inv_1 U257 (.A(n160), .Y(n194));
sg13g2_inv_1 U258 (.A(n158), .Y(n198));
sg13g2_inv_1 U259 (.A(n155), .Y(n195));
sg13g2_inv_1 U260 (.A(n162), .Y(n197));
sg13g2_xor2_1 U261 (.A(N13), .B(n217), .X(N727));
sg13g2_nor2_1 U262 (.A(n190), .B(n218), .Y(n217));
sg13g2_xor2_1 U263 (.A(N9), .B(n219), .X(N726));
sg13g2_nor2_1 U264 (.A(n165), .B(n218), .Y(n219));
sg13g2_xor2_1 U265 (.A(N5), .B(n220), .X(N725));
sg13g2_nor2_1 U266 (.A(n188), .B(n218), .Y(n220));
sg13g2_xor2_1 U267 (.A(N1), .B(n221), .X(N724));
sg13g2_nor2_1 U268 (.A(n163), .B(n218), .Y(n221));
sg13g2_nand4_1 U269 (.A(n155), .B(n193), .C(n160), .D(n204), .Y(n218));
sg13g2_nand2_1 U270 (.A(n222), .B(n223), .Y(n204));
sg13g2_or3_1 U271 (.A(n189), .B(n176), .C(n172), .X(n223));
sg13g2_inv_1 U272 (.A(n188), .Y(n172));
sg13g2_inv_1 U273 (.A(n190), .Y(n176));
sg13g2_nor2_1 U274 (.A(n165), .B(n163), .Y(n189));
sg13g2_or3_1 U275 (.A(n164), .B(n173), .C(n175), .X(n222));
sg13g2_inv_1 U276 (.A(n163), .Y(n175));
sg13g2_inv_1 U277 (.A(n165), .Y(n173));
sg13g2_xor2_1 U278 (.A(n224), .B(n225), .X(n165));
sg13g2_xor2_1 U279 (.A(n226), .B(n227), .X(n225));
sg13g2_xor2_1 U280 (.A(N25), .B(N105), .X(n227));
sg13g2_xor2_1 U281 (.A(N97), .B(N9), .X(n226));
sg13g2_xor2_1 U282 (.A(n228), .B(n229), .X(n224));
sg13g2_xor2_1 U283 (.A(n230), .B(n231), .X(n229));
sg13g2_xor2_1 U284 (.A(n232), .B(n233), .X(n228));
sg13g2_nand2_1 U285 (.A(N131), .B(N137), .Y(n232));
sg13g2_nor2_1 U286 (.A(n190), .B(n188), .Y(n164));
sg13g2_xor2_1 U287 (.A(n234), .B(n235), .X(n188));
sg13g2_xor2_1 U288 (.A(n236), .B(n237), .X(n234));
sg13g2_xor2_1 U289 (.A(n238), .B(n239), .X(n237));
sg13g2_xor2_1 U290 (.A(N121), .B(N109), .X(n239));
sg13g2_xor2_1 U291 (.A(N21), .B(N125), .X(n238));
sg13g2_xor2_1 U292 (.A(n240), .B(n241), .X(n236));
sg13g2_xor2_1 U293 (.A(n242), .B(n243), .X(n241));
sg13g2_xor2_1 U294 (.A(n244), .B(N101), .X(n240));
sg13g2_nand2_1 U295 (.A(N130), .B(N137), .Y(n244));
sg13g2_xor2_1 U296 (.A(n245), .B(n246), .X(n190));
sg13g2_xor2_1 U297 (.A(n247), .B(n248), .X(n246));
sg13g2_xor2_1 U298 (.A(N117), .B(N113), .X(n248));
sg13g2_xor2_1 U299 (.A(N81), .B(N13), .X(n247));
sg13g2_xor2_1 U300 (.A(n249), .B(n250), .X(n245));
sg13g2_xor2_1 U301 (.A(n251), .B(n252), .X(n250));
sg13g2_nand2_1 U302 (.A(N132), .B(N137), .Y(n251));
sg13g2_xor2_1 U303 (.A(n253), .B(n254), .X(n249));
sg13g2_xor2_1 U304 (.A(n255), .B(n256), .X(n160));
sg13g2_xor2_1 U305 (.A(n235), .B(n257), .X(n256));
sg13g2_xor2_1 U306 (.A(n258), .B(n259), .X(n257));
sg13g2_nand2_1 U307 (.A(N134), .B(N137), .Y(n259));
sg13g2_inv_1 U308 (.A(N57), .Y(n258));
sg13g2_xor2_1 U309 (.A(N117), .B(n260), .X(n235));
sg13g2_xor2_1 U310 (.A(N53), .B(N37), .X(n260));
sg13g2_xor2_1 U311 (.A(n261), .B(n230), .X(n255));
sg13g2_xor2_1 U312 (.A(N101), .B(n262), .X(n230));
sg13g2_xor2_1 U313 (.A(N69), .B(N41), .X(n262));
sg13g2_xor2_1 U314 (.A(n253), .B(n263), .X(n261));
sg13g2_xnor2_1 U315 (.A(N45), .B(n264), .Y(n253));
sg13g2_xor2_1 U316 (.A(N85), .B(N61), .X(n264));
sg13g2_nor2_1 U317 (.A(n162), .B(n158), .Y(n193));
sg13g2_xor2_1 U318 (.A(n265), .B(n266), .X(n158));
sg13g2_xor2_1 U319 (.A(N73), .B(N33), .X(n266));
sg13g2_xor2_1 U320 (.A(n267), .B(n268), .X(n265));
sg13g2_xor2_1 U321 (.A(n269), .B(n270), .X(n268));
sg13g2_xor2_1 U322 (.A(N37), .B(N1), .X(n270));
sg13g2_xor2_1 U323 (.A(N45), .B(N41), .X(n269));
sg13g2_xor2_1 U324 (.A(n271), .B(n272), .X(n267));
sg13g2_xor2_1 U325 (.A(n254), .B(n273), .X(n272));
sg13g2_xor2_1 U326 (.A(N121), .B(N89), .X(n254));
sg13g2_xor2_1 U327 (.A(n274), .B(n242), .X(n271));
sg13g2_xor2_1 U328 (.A(N105), .B(N5), .X(n242));
sg13g2_nand2_1 U329 (.A(N137), .B(N135), .Y(n274));
sg13g2_xor2_1 U330 (.A(n275), .B(n276), .X(n162));
sg13g2_xor2_1 U331 (.A(n277), .B(n278), .X(n276));
sg13g2_xor2_1 U332 (.A(n279), .B(n280), .X(n278));
sg13g2_nand2_1 U333 (.A(N133), .B(N137), .Y(n280));
sg13g2_inv_1 U334 (.A(N29), .Y(n279));
sg13g2_xor2_1 U335 (.A(N65), .B(N5), .X(n277));
sg13g2_xor2_1 U336 (.A(n281), .B(n282), .X(n275));
sg13g2_xor2_1 U337 (.A(n283), .B(n273), .X(n282));
sg13g2_xor2_1 U338 (.A(N13), .B(N9), .X(n273));
sg13g2_xor2_1 U339 (.A(n284), .B(n243), .X(n281));
sg13g2_xor2_1 U340 (.A(N113), .B(N97), .X(n243));
sg13g2_xor2_1 U341 (.A(n285), .B(n286), .X(n155));
sg13g2_xor2_1 U342 (.A(n287), .B(n288), .X(n286));
sg13g2_xor2_1 U343 (.A(N49), .B(N17), .X(n288));
sg13g2_xor2_1 U344 (.A(N61), .B(N53), .X(n287));
sg13g2_xor2_1 U345 (.A(n289), .B(n290), .X(n285));
sg13g2_xor2_1 U346 (.A(n291), .B(n252), .X(n290));
sg13g2_xnor2_1 U347 (.A(N125), .B(n292), .Y(n252));
sg13g2_xor2_1 U348 (.A(N93), .B(N29), .X(n292));
sg13g2_nand2_1 U349 (.A(N136), .B(N137), .Y(n291));
sg13g2_xnor2_1 U350 (.A(n233), .B(n283), .Y(n289));
sg13g2_xor2_1 U351 (.A(N21), .B(N25), .X(n283));
sg13g2_xor2_1 U352 (.A(N109), .B(n293), .X(n233));
sg13g2_xor2_1 U353 (.A(N77), .B(N57), .X(n293));
sg13g2_xor2_1 U354 (.A(n294), .B(N85), .X(n163));
sg13g2_xor2_1 U355 (.A(n295), .B(n296), .X(n294));
sg13g2_xor2_1 U356 (.A(n297), .B(n298), .X(n296));
sg13g2_xor2_1 U357 (.A(N77), .B(N69), .X(n298));
sg13g2_xor2_1 U358 (.A(N93), .B(N89), .X(n297));
sg13g2_xor2_1 U359 (.A(n299), .B(n300), .X(n295));
sg13g2_xor2_1 U360 (.A(n263), .B(n231), .X(n300));
sg13g2_xor2_1 U361 (.A(N65), .B(N73), .X(n231));
sg13g2_xor2_1 U362 (.A(N33), .B(N49), .X(n263));
sg13g2_xor2_1 U363 (.A(n301), .B(n302), .X(n299));
sg13g2_inv_1 U364 (.A(n284), .Y(n302));
sg13g2_xnor2_1 U365 (.A(N1), .B(n303), .Y(n284));
sg13g2_xor2_1 U366 (.A(N81), .B(N17), .X(n303));
sg13g2_nand2_1 U367 (.A(N129), .B(N137), .Y(n301));
endmodule

